



<!DOCTYPE html>
<html lang="es-SV">

<head>
<title>Directorio de empresas de El Salvador | P&aacute;ginas Amarillas</title>
<link rel="canonical" href="http://www.paginasamarillas.com.sv" />
<meta name="description"
	content="P&aacute;ginas Amarillas de Publicar es el directorio m&aacute;s completo de El Salvador. En nuestra gu&iacute;a de empresas podr&aacute; solicitar toda la informaci&oacute;n comercial de empresas, productos y servicios en El Salvador.">


<!--head-->




<!-- Google Tag Manager -->
<noscript>
	<iframe
		src="//www.googletagmanager.com/ns.html?id=GTM-WTPB5H"
		height="0" width="0" style="display:none;visibility:hidden"></iframe>
</noscript>
<script>
	(function(w, d, s, l, i) {
		w[l] = w[l] || [];
		w[l].push({
			'gtm.start' : new Date().getTime(),
			event : 'gtm.js'
		});
		var f = d.getElementsByTagName(s)[0], j = d.createElement(s), dl = l != 'dataLayer' ? '&l='
				+ l
				: '';
		j.async = true;
		j.src = '//www.googletagmanager.com/gtm.js?id=' + i + dl;
		f.parentNode.insertBefore(j, f);
	})(window, document, 'script', 'dataLayer',
			'GTM-WTPB5H');
</script>
<!-- End Google Tag Manager -->

<meta charset="UTF-8">
<meta http-equiv="X-UA-Compatible" content="IE=edge">
<!-- <meta name="viewport" content="width=device-width, initial-scale=1"> -->
<meta name="viewport" content="width=1024">

<!-- Meta SuTarget Publisher -->

<meta name="cXenseParse:publishername" content="PAGINASMARILLAS">
<meta name="cXenseParse:pageclass" content="frontpage">
<meta name="cXenseParse:recs:recommendable" content="false">
<!-- End Meta SuTarget Publisher -->

<link rel="shortcut icon" href="/view/global/common/images/favicon.ico" type="image/x-icon" />

<!--Reset-->
<link href="/view/global/common/css/normalize.css" rel="stylesheet">
<!-- Bootstrap -->
<link href="/view/global/common/vendor/bootstrap/css/bootstrap.min.css" rel="stylesheet">
<!--estilos fuentes-->
<link href="/view/global/common/css/fonts.css?20171115" rel="stylesheet">
<!--estilos main-->
<link href="/view/global/common/css/main.css?20171207" rel="stylesheet">

<!--Comienzo de llamados necesarios para analytics -->
<script src="/view/global/common/vendor/jquery/jquery-3.2.1.min.js"></script>
<script src="/view/global/common/js/sessionStorage_utils.js"></script>
<script type="text/javascript">
	var directoryIdJsp = "1";
</script>





   
      
   
        
   		<script type="text/javascript">
	var HAF = {};
	HAF.config = {'global':{'internalDomains':'javascript:,ar.amarillas.dev.yellargentina.com','trackDownloadLinks':true,'charset':'UTF-8','trackExternalLinks':false,'currenty':'ARS','fwjsurl':'/view/common/js/analytics/yell-analytics.js?20170630'},'stc':{'server':'http://dzmkkiowi0jbc.cloudfront.net','country':2,'url.path':'/js/las/analytics.js','account':1111,'enabled':true}}
</script>
<script type="text/javascript" charset="UTF-8" src="http://dzmkkiowi0jbc.cloudfront.net/js/las/analytics.js"></script>
<script type="text/javascript" charset="UTF-8" src="/view/common/js/analytics/yell-analytics.js?20170630"></script>

   
   
   
    
   
   
    
   



<!--Final de llamados necesarios para analytics -->

<!-- HTML5 shim and Respond.js for IE8 support of HTML5 elements and media queries -->
<!-- WARNING: Respond.js doesn't work if you view the page via file:// -->
<!--[if lt IE 9]>
  <script src="https://oss.maxcdn.com/html5shiv/3.7.3/html5shiv.min.js"></script>
  <script src="https://oss.maxcdn.com/respond/1.4.2/respond.min.js"></script>
<![endif]-->



	
	


<!--URL Independientes-->
<!--<link media="media=only screen and (max-width: 640px)" href="http://m.paginasamarillas.com.sv/" />-->




<!-- Cxense script start -->
<script id="navegg" type="text/javascript" src="//tag.navdmp.com/tm21360.js"></script>
<script type="text/javascript">
nvg21360.makeCustomSegment = function (){ var res = {}; this.cokCache = {}; var nvg_parms = new Array('gender', 'age', 'education', 'interest', 'product', 'income', 'marital', 'prolook'); for (nvg_i in nvg_parms) { var nvg_tmp_arr = ''; var nvg_tmp_nme = nvg_parms[nvg_i]; var nvg_tmp = this.getSegment(nvg_parms[nvg_i]); if (nvg_tmp.search(',') != -1) { res[ nvg_tmp_nme ] = nvg_tmp.split(','); } else if (nvg_tmp.search('-') != -1) { res[ nvg_tmp_nme ] = nvg_tmp.split('-'); } else if (nvg_tmp != '') { res[ nvg_tmp_nme ] = nvg_tmp; } } return res; };
const segments = nvg21360.makeCustomSegment();
</script>
<script>
var cX = cX || {}; cX.callQueue = cX.callQueue || [];
cX.callQueue.push(['setSiteId', '1129412760827754572']);
cX.callQueue.push(['setUserProfileParameters', segments ]);
cX.callQueue.push(['sendPageViewEvent']);
</script>
<script type="text/javascript">
(function(d,s,e,t){e=d.createElement(s);e.type='text/java'+s;e.async='async';
e.src='http'+('https:'===location.protocol?'s://s':'://')+'cdn.cxense.com/cx.js';
t=d.getElementsByTagName(s)[0];t.parentNode.insertBefore(e,t);})(document,'script');
</script>
<!-- Cxense script end -->


	<!-- Start Alexa Certify Javascript -->
	<script type="text/javascript">
	_atrk_opts = { atrk_acct:"m480m1aQibl0T3", domain:"paginasamarillas.com.sv",dynamic: true};
	(function() { var as = document.createElement('script'); as.type = 'text/javascript'; as.async = true; as.src = "https://d31qbv1cthcecs.cloudfront.net/atrk.js"; var s = document.getElementsByTagName('script')[0];s.parentNode.insertBefore(as, s); })();
	</script>
	<noscript><img src="https://d5nxst8fruw4z.cloudfront.net/atrk.gif?account=m480m1aQibl0T3" style="display:none" height="1" width="1" alt="" /></noscript>
	<!-- End Alexa Certify Javascript -->


<!-- Facebook Pixel Code -->
<script>
  !function(f,b,e,v,n,t,s)
  {if(f.fbq)return;n=f.fbq=function(){n.callMethod?
  n.callMethod.apply(n,arguments):n.queue.push(arguments)};
  if(!f._fbq)f._fbq=n;n.push=n;n.loaded=!0;n.version='2.0';
  n.queue=[];t=b.createElement(e);t.async=!0;
  t.src=v;s=b.getElementsByTagName(e)[0];
  s.parentNode.insertBefore(t,s)}(window, document,'script',
  'https://connect.facebook.net/en_US/fbevents.js');
  fbq('init', '147004932590647');
  fbq('track', 'PageView');
</script>
<noscript><img height="1" width="1" style="display:none"
  src="https://www.facebook.com/tr?id=147004932590647&ev=PageView&noscript=1"
/></noscript>
<!-- End Facebook Pixel Code -->

<!--home main-->
<link href="/view/global/common/css/home.css?20170906" rel="stylesheet">


 <!-- Start Alexa Certify Javascript -->
 <script type="text/javascript"> _atrk_opts = { atrk_acct:"m480m1aQibl0T3", domain:"paginasamarillas.com.sv",dynamic: true}; (function() { var as = document.createElement('script'); as.type = 'text/javascript'; as.async = true; as.src = "https://d31qbv1cthcecs.cloudfront.net/atrk.js"; var s = document.getElementsByTagName('script')[0];s.parentNode.insertBefore(as, s); })();</script> 
 
 <noscript><img src="https://d5nxst8fruw4z.cloudfront.net/atrk.gif?account=m480m1aQibl0T3" style="display:none" height="1" width="1" alt="" /></noscript><!-- End Alexa Certify Javascript --> 


 
<style>
.homeBg {
	background-image:
		url(/view/global/common/images/backgrounds/6.jpg);
}
</style>
</head>

<body class="home">
	

<!-- Google Tag Manager (noscript) -->
<noscript><iframe src="https://www.googletagmanager.com/ns.html?id=GTM-WTPB5H" height="0" width="0" style="display:none;visibility:hidden"></iframe></noscript>
<!-- End Google Tag Manager (noscript) -->

	<section class="main">
		<!--fixed top menu-->
		



<header class="top">
    <div class="container">
        <div class="top-left">
            <ul class="top-list">
                <a href="/">
                    <i class="pa-icon logo-small"></i>
                </a>
            </ul>
		</div>
		<div class="top-center">
			<div class="logoHome pa-icon"></div>
			<div class="search">
				<h1 class="">Páginas amarillas de
					<span class="countryTitle">El Salvador</span>
				</h1>
				<div class="homeTxt">El directorio más completo de <strong>Latinoamérica</strong> a un clic de distancia</div>
			</div>

			<form id="searchForm" class="formCity search-form" role="search">
				<div class="searchContain">
					<div class="elementForm">
						<input id="keyword" data-container="body" data-toggle="popover" data-placement="bottom" data-content="Ingrese al menos 2 caracteres" type="text" class="form-control what-field" value="" placeholder="&iquest;Qu&eacute; buscas&#63;" autocomplete="off">
					</div>
					<div class="elementForm">
						<input id="locality" type="text" class="form-control where-field" value="" placeholder="&iquest;D&oacute;nde&#63;" autocomplete="off">
					</div>
					<input type="hidden" id="friendlyName" name="friendlyName">
					<button id="buscar" type="submit" class="btn btn-default icon-pa_02 searchSite" disabled></button>
				</div>

				<div class="m-suggest hide" id="suggestions">
					<span class="suggarrow-shadow"></span><span class="suggarrow"></span>
					<div></div>
				</div>
				<div class="m-suggest hide" id="suggestionsLocality">
					<span class="suggarrow-shadow"></span><span class="suggarrow"></span>
					<div></div>
				</div>
			</form>
			
			
            
		</div>
		<div class="top-right">
			<ul class="top-list">
				<li>
					<span class="icon-pa_03"></span>
					<span class="is-link topButton" data-toggle="modal" data-target="#anuncia-modal" target="_blank" title="Anuncia con nosotros">Anúnciate</span>
                </li>
                
	                <li class="printGuide">
						<span class="icon-pa_66"></span>
						<a class="is-link topButton" href="http://sites.paginasamarillas.com/directorio/home.html" target="_blank" onclick="return clickGuidePrinted(this,TipoClick.CLIC_WEB,Pagina.PAGE_HOME);">Guía Impresa</a>
	                </li>
                
                <li>
                   <!--seleccionar ciudad popover-->
                   <div class="countrySelect">
                       <span class="icon-pa_04"></span>
                       

	                       <div class="topButton " data-popover="placeSelect" id="place" data-placement="bottom" data-popover-fixed data-toggle="popover" data-container="body" data-html="true">
	                       		<div class="citynameWrap">
	                       			El Salvador
	                       		</div>
	                       	<span class=" drop icon-pa_01 "></span> 
	                       </div>
                       
              
                       
                       <div id="placeSelect" class="hide popover-custom center">
                           <form class="dataForm countryForm form-inline" role="form" action="/" method="post">
                               <div class="row">
                                   <div class="form-group col-xs-12">
                                        <label for="search-countrySelect" class="bold control-label selectTitle">&iquest;En qué país te encuentras&#63;</label>
	                                    <div class="selectWrap">
	                                        <select id="search-countrySelect" class="form-control input-sm regular search-countrySelect">
	                                        	

	                                        	
	                                        		<option value="http://www.paginasamarillas.com.ar/" >Argentina</option>
	                                        	
	                                        		<option value="http://bolivia.paginasamarillas.com/" >Bolivia</option>
	                                        	
	                                        		<option value="http://www.amarillas.cl/ " >Chile</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.co/" >Colombia</option>
	                                        	
	                                        		<option value="http://costa-rica.paginasamarillas.com/" >Costa Rica</option>
	                                        	
	                                        		<option value="http://www.paginas-amarillas.com.ec/" >Ecuador</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.sv/" selected>El Salvador</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.gt/" >Guatemala</option>
	                                        	
	                                        		<option value="http://honduras.paginasamarillas.com/" >Honduras</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com/latinoamerica" >Latinoamerica</option>
	                                        	
	                                        		<option value="http://mexico.paginasamarillas.com/" >Mexico</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.ni/" >Nicaragua</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.pa/" >Panamá</option>
	                                        	
	                                        		<option value="http://www.paginasamarillas.com.pe/" >Perú</option>
	                                        	
	                                        		<option value="http://puerto-rico.paginasamarillas.com/" >Puerto Rico</option>
	                                        	
	                                        		<option value="http://republica-dominicana.paginasamarillas.com/" >República Dominicana</option>
	                                        	
	                                        		<option value="http://venezuela.paginasamarillas.com/" >Venezuela</option>
	                                        	
	                                        </select>
	                                        <button type="submit" class="btn btnGps blueBtn icon-pa_33 city"></button>
	                                    </div>
                                	</div>

									<div class="form-group col-xs-12">
										<label for="search-citySelect" class="bold control-label selectTitle">&iquest;En qué ciudad&#63;</label>
										<div class="selectWrap">
											<select id="search-citySelect" class="form-control input-sm regular search-citySelect" name="city-selector">
												<option value="">Todas las ciudades</option>
		                                        
		                                        	
	                                        	
		                                        	
		                                        		<option value="Cochabamba"
		                                        			class="hide c1"
		                                        			>Cochabamba</option>
		                                        	
		                                        		<option value="Chuquisaca"
		                                        			class="hide c1"
		                                        			>Chuquisaca</option>
		                                        	
		                                        		<option value="El Alto"
		                                        			class="hide c1"
		                                        			>El Alto</option>
		                                        	
		                                        		<option value="Montero"
		                                        			class="hide c1"
		                                        			>Montero</option>
		                                        	
		                                        		<option value="La Paz"
		                                        			class="hide c1"
		                                        			>La Paz</option>
		                                        	
		                                        		<option value="Potosi"
		                                        			class="hide c1"
		                                        			>Potosi</option>
		                                        	
		                                        		<option value="Oruro"
		                                        			class="hide c1"
		                                        			>Oruro</option>
		                                        	
		                                        		<option value="Santa Cruz"
		                                        			class="hide c1"
		                                        			>Santa Cruz</option>
		                                        	
		                                        		<option value="Sucre"
		                                        			class="hide c1"
		                                        			>Sucre</option>
		                                        	
		                                        		<option value="Tarija"
		                                        			class="hide c1"
		                                        			>Tarija</option>
		                                        	
		                                        		<option value="Urbana"
		                                        			class="hide c1"
		                                        			>Urbana</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Santiago de Chile"
		                                        			class="hide c2"
		                                        			>Santiago de Chile</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Bogotá"
		                                        			class="hide c3"
		                                        			>Bogotá</option>
		                                        	
		                                        		<option value="Medellín"
		                                        			class="hide c3"
		                                        			>Medellín</option>
		                                        	
		                                        		<option value="Cali"
		                                        			class="hide c3"
		                                        			>Cali</option>
		                                        	
		                                        		<option value="Barranquilla"
		                                        			class="hide c3"
		                                        			>Barranquilla</option>
		                                        	
		                                        		<option value="Cartagena de Indias"
		                                        			class="hide c3"
		                                        			>Cartagena de Indias</option>
		                                        	
		                                        		<option value="Cúcuta"
		                                        			class="hide c3"
		                                        			>Cúcuta</option>
		                                        	
		                                        		<option value="Ibague"
		                                        			class="hide c3"
		                                        			>Ibague</option>
		                                        	
		                                        		<option value="Bucaramanga"
		                                        			class="hide c3"
		                                        			>Bucaramanga</option>
		                                        	
		                                        		<option value="Santa Marta"
		                                        			class="hide c3"
		                                        			>Santa Marta</option>
		                                        	
		                                        		<option value="Villavicencio"
		                                        			class="hide c3"
		                                        			>Villavicencio</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Alajuela"
		                                        			class="hide c4"
		                                        			>Alajuela</option>
		                                        	
		                                        		<option value="Barva"
		                                        			class="hide c4"
		                                        			>Barva</option>
		                                        	
		                                        		<option value="Cartago"
		                                        			class="hide c4"
		                                        			>Cartago</option>
		                                        	
		                                        		<option value="Guadalupe"
		                                        			class="hide c4"
		                                        			>Guadalupe</option>
		                                        	
		                                        		<option value="Guanacaste"
		                                        			class="hide c4"
		                                        			>Guanacaste</option>
		                                        	
		                                        		<option value="Heredia"
		                                        			class="hide c4"
		                                        			>Heredia</option>
		                                        	
		                                        		<option value="Liberia"
		                                        			class="hide c4"
		                                        			>Liberia</option>
		                                        	
		                                        		<option value="Limón"
		                                        			class="hide c4"
		                                        			>Limón</option>
		                                        	
		                                        		<option value="Puntaresnas"
		                                        			class="hide c4"
		                                        			>Puntaresnas</option>
		                                        	
		                                        		<option value="San José"
		                                        			class="hide c4"
		                                        			>San José</option>
		                                        	
		                                        		<option value="Uruca"
		                                        			class="hide c4"
		                                        			>Uruca</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Ambato"
		                                        			class="hide c5"
		                                        			>Ambato</option>
		                                        	
		                                        		<option value="Cuenca"
		                                        			class="hide c5"
		                                        			>Cuenca</option>
		                                        	
		                                        		<option value="Durán"
		                                        			class="hide c5"
		                                        			>Durán</option>
		                                        	
		                                        		<option value="Guayaquil"
		                                        			class="hide c5"
		                                        			>Guayaquil</option>
		                                        	
		                                        		<option value="Manta"
		                                        			class="hide c5"
		                                        			>Manta</option>
		                                        	
		                                        		<option value="Machala"
		                                        			class="hide c5"
		                                        			>Machala</option>
		                                        	
		                                        		<option value="Portoviejo"
		                                        			class="hide c5"
		                                        			>Portoviejo</option>
		                                        	
		                                        		<option value="Loja"
		                                        			class="hide c5"
		                                        			>Loja</option>
		                                        	
		                                        		<option value="Quito"
		                                        			class="hide c5"
		                                        			>Quito</option>
		                                        	
		                                        		<option value="Santo Domingo"
		                                        			class="hide c5"
		                                        			>Santo Domingo</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Ahuachapán"
		                                        			class=" c6"
		                                        			>Ahuachapán</option>
		                                        	
		                                        		<option value="Chalatenango"
		                                        			class=" c6"
		                                        			>Chalatenango</option>
		                                        	
		                                        		<option value="Cojutepeque"
		                                        			class=" c6"
		                                        			>Cojutepeque</option>
		                                        	
		                                        		<option value="La Unión"
		                                        			class=" c6"
		                                        			>La Unión</option>
		                                        	
		                                        		<option value="Santa Ana"
		                                        			class=" c6"
		                                        			>Santa Ana</option>
		                                        	
		                                        		<option value="San Francisco Gotera"
		                                        			class=" c6"
		                                        			>San Francisco Gotera</option>
		                                        	
		                                        		<option value="San Miguel"
		                                        			class=" c6"
		                                        			>San Miguel</option>
		                                        	
		                                        		<option value="San Salvador"
		                                        			class=" c6"
		                                        			>San Salvador</option>
		                                        	
		                                        		<option value="San Vicente"
		                                        			class=" c6"
		                                        			>San Vicente</option>
		                                        	
		                                        		<option value="Sensuntepeque"
		                                        			class=" c6"
		                                        			>Sensuntepeque</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Huehuetenango "
		                                        			class="hide c7"
		                                        			>Huehuetenango </option>
		                                        	
		                                        		<option value="Santa Cruz del Quiché "
		                                        			class="hide c7"
		                                        			>Santa Cruz del Quiché </option>
		                                        	
		                                        		<option value="Chimaltenango "
		                                        			class="hide c7"
		                                        			>Chimaltenango </option>
		                                        	
		                                        		<option value="Guatemala "
		                                        			class="hide c7"
		                                        			>Guatemala </option>
		                                        	
		                                        		<option value="Coban "
		                                        			class="hide c7"
		                                        			>Coban </option>
		                                        	
		                                        		<option value="Escuintla "
		                                        			class="hide c7"
		                                        			>Escuintla </option>
		                                        	
		                                        		<option value="Mazatenango "
		                                        			class="hide c7"
		                                        			>Mazatenango </option>
		                                        	
		                                        		<option value="Quetzaltenango "
		                                        			class="hide c7"
		                                        			>Quetzaltenango </option>
		                                        	
		                                        		<option value="Flores "
		                                        			class="hide c7"
		                                        			>Flores </option>
		                                        	
		                                        		<option value="San Marcos "
		                                        			class="hide c7"
		                                        			>San Marcos </option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Tegucigalpa"
		                                        			class="hide c8"
		                                        			>Tegucigalpa</option>
		                                        	
		                                        		<option value="San Pedro Sula"
		                                        			class="hide c8"
		                                        			>San Pedro Sula</option>
		                                        	
		                                        		<option value="La Ceiba"
		                                        			class="hide c8"
		                                        			>La Ceiba</option>
		                                        	
		                                        		<option value="Choloma"
		                                        			class="hide c8"
		                                        			>Choloma</option>
		                                        	
		                                        		<option value="Danlí"
		                                        			class="hide c8"
		                                        			>Danlí</option>
		                                        	
		                                        		<option value="Choluteca"
		                                        			class="hide c8"
		                                        			>Choluteca</option>
		                                        	
		                                        		<option value="Juticalpa"
		                                        			class="hide c8"
		                                        			>Juticalpa</option>
		                                        	
		                                        		<option value="Catacamas"
		                                        			class="hide c8"
		                                        			>Catacamas</option>
		                                        	
		                                        		<option value="Comayagua"
		                                        			class="hide c8"
		                                        			>Comayagua</option>
		                                        	
		                                        		<option value="Santa Rosa De Copán"
		                                        			class="hide c8"
		                                        			>Santa Rosa De Copán</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Bogotá"
		                                        			class="hide c9"
		                                        			>Bogotá</option>
		                                        	
		                                        		<option value="La Paz"
		                                        			class="hide c9"
		                                        			>La Paz</option>
		                                        	
		                                        		<option value="Santiago de Chile"
		                                        			class="hide c9"
		                                        			>Santiago de Chile</option>
		                                        	
		                                        		<option value="San José"
		                                        			class="hide c9"
		                                        			>San José</option>
		                                        	
		                                        		<option value="Quito"
		                                        			class="hide c9"
		                                        			>Quito</option>
		                                        	
		                                        		<option value="San Salvador"
		                                        			class="hide c9"
		                                        			>San Salvador</option>
		                                        	
		                                        		<option value="Ciudad de Guatemala"
		                                        			class="hide c9"
		                                        			>Ciudad de Guatemala</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Baja California"
		                                        			class="hide c10"
		                                        			>Baja California</option>
		                                        	
		                                        		<option value="Baja California Sur"
		                                        			class="hide c10"
		                                        			>Baja California Sur</option>
		                                        	
		                                        		<option value="Campeche"
		                                        			class="hide c10"
		                                        			>Campeche</option>
		                                        	
		                                        		<option value="Chiapas"
		                                        			class="hide c10"
		                                        			>Chiapas</option>
		                                        	
		                                        		<option value="Chihuahua"
		                                        			class="hide c10"
		                                        			>Chihuahua</option>
		                                        	
		                                        		<option value="Colima"
		                                        			class="hide c10"
		                                        			>Colima</option>
		                                        	
		                                        		<option value="Jalisco"
		                                        			class="hide c10"
		                                        			>Jalisco</option>
		                                        	
		                                        		<option value="Mexico"
		                                        			class="hide c10"
		                                        			>Mexico</option>
		                                        	
		                                        		<option value="Morellia"
		                                        			class="hide c10"
		                                        			>Morellia</option>
		                                        	
		                                        		<option value="Puebla"
		                                        			class="hide c10"
		                                        			>Puebla</option>
		                                        	
		                                        		<option value="Tabasco"
		                                        			class="hide c10"
		                                        			>Tabasco</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Matagalpa"
		                                        			class="hide c11"
		                                        			>Matagalpa</option>
		                                        	
		                                        		<option value="Chinandega"
		                                        			class="hide c11"
		                                        			>Chinandega</option>
		                                        	
		                                        		<option value="Estelí"
		                                        			class="hide c11"
		                                        			>Estelí</option>
		                                        	
		                                        		<option value="Granada"
		                                        			class="hide c11"
		                                        			>Granada</option>
		                                        	
		                                        		<option value="Ciudad Sandino"
		                                        			class="hide c11"
		                                        			>Ciudad Sandino</option>
		                                        	
		                                        		<option value="León"
		                                        			class="hide c11"
		                                        			>León</option>
		                                        	
		                                        		<option value="Managua"
		                                        			class="hide c11"
		                                        			>Managua</option>
		                                        	
		                                        		<option value="Masaya"
		                                        			class="hide c11"
		                                        			>Masaya</option>
		                                        	
		                                        		<option value="Juigalpa"
		                                        			class="hide c11"
		                                        			>Juigalpa</option>
		                                        	
		                                        		<option value="Tipitapa"
		                                        			class="hide c11"
		                                        			>Tipitapa</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Panamá"
		                                        			class="hide c12"
		                                        			>Panamá</option>
		                                        	
		                                        		<option value="David"
		                                        			class="hide c12"
		                                        			>David</option>
		                                        	
		                                        		<option value="Colón"
		                                        			class="hide c12"
		                                        			>Colón</option>
		                                        	
		                                        		<option value="Penonomé"
		                                        			class="hide c12"
		                                        			>Penonomé</option>
		                                        	
		                                        		<option value="Santiago"
		                                        			class="hide c12"
		                                        			>Santiago</option>
		                                        	
		                                        		<option value="Bocas del Toro"
		                                        			class="hide c12"
		                                        			>Bocas del Toro</option>
		                                        	
		                                        		<option value="Chitré"
		                                        			class="hide c12"
		                                        			>Chitré</option>
		                                        	
		                                        		<option value="Las Tablas"
		                                        			class="hide c12"
		                                        			>Las Tablas</option>
		                                        	
		                                        		<option value="Las Palmas"
		                                        			class="hide c12"
		                                        			>Las Palmas</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Arequipa"
		                                        			class="hide c13"
		                                        			>Arequipa</option>
		                                        	
		                                        		<option value="Ayacucho"
		                                        			class="hide c13"
		                                        			>Ayacucho</option>
		                                        	
		                                        		<option value="Cuzco"
		                                        			class="hide c13"
		                                        			>Cuzco</option>
		                                        	
		                                        		<option value="Huanuco"
		                                        			class="hide c13"
		                                        			>Huanuco</option>
		                                        	
		                                        		<option value="Ica"
		                                        			class="hide c13"
		                                        			>Ica</option>
		                                        	
		                                        		<option value="Junin"
		                                        			class="hide c13"
		                                        			>Junin</option>
		                                        	
		                                        		<option value="Lima"
		                                        			class="hide c13"
		                                        			>Lima</option>
		                                        	
		                                        		<option value="Esqui"
		                                        			class="hide c13"
		                                        			>Esqui</option>
		                                        	
		                                        		<option value="Pasco"
		                                        			class="hide c13"
		                                        			>Pasco</option>
		                                        	
		                                        		<option value="Piura"
		                                        			class="hide c13"
		                                        			>Piura</option>
		                                        	
		                                        		<option value="Tumbes"
		                                        			class="hide c13"
		                                        			>Tumbes</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Altamira"
		                                        			class="hide c14"
		                                        			>Altamira</option>
		                                        	
		                                        		<option value="Arecibo"
		                                        			class="hide c14"
		                                        			>Arecibo</option>
		                                        	
		                                        		<option value="Bayamón"
		                                        			class="hide c14"
		                                        			>Bayamón</option>
		                                        	
		                                        		<option value="Barranquitas"
		                                        			class="hide c14"
		                                        			>Barranquitas</option>
		                                        	
		                                        		<option value="Carolina"
		                                        			class="hide c14"
		                                        			>Carolina</option>
		                                        	
		                                        		<option value="Humacao"
		                                        			class="hide c14"
		                                        			>Humacao</option>
		                                        	
		                                        		<option value="Guayama"
		                                        			class="hide c14"
		                                        			>Guayama</option>
		                                        	
		                                        		<option value="Mayagues"
		                                        			class="hide c14"
		                                        			>Mayagues</option>
		                                        	
		                                        		<option value="Ponce"
		                                        			class="hide c14"
		                                        			>Ponce</option>
		                                        	
		                                        		<option value="Puerto Rico"
		                                        			class="hide c14"
		                                        			>Puerto Rico</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Cibao"
		                                        			class="hide c15"
		                                        			>Cibao</option>
		                                        	
		                                        		<option value="Baoruco"
		                                        			class="hide c15"
		                                        			>Baoruco</option>
		                                        	
		                                        		<option value="Duarte"
		                                        			class="hide c15"
		                                        			>Duarte</option>
		                                        	
		                                        		<option value="Espaillat"
		                                        			class="hide c15"
		                                        			>Espaillat</option>
		                                        	
		                                        		<option value="Higuet"
		                                        			class="hide c15"
		                                        			>Higuet</option>
		                                        	
		                                        		<option value="La Vega"
		                                        			class="hide c15"
		                                        			>La Vega</option>
		                                        	
		                                        		<option value="La Romana"
		                                        			class="hide c15"
		                                        			>La Romana</option>
		                                        	
		                                        		<option value="Puerto Plata"
		                                        			class="hide c15"
		                                        			>Puerto Plata</option>
		                                        	
		                                        		<option value="Santiago"
		                                        			class="hide c15"
		                                        			>Santiago</option>
		                                        	
		                                        		<option value="Santo Domingo"
		                                        			class="hide c15"
		                                        			>Santo Domingo</option>
		                                        	
		                                        		<option value="Samana"
		                                        			class="hide c15"
		                                        			>Samana</option>
		                                        	
	                                        	
		                                        	
		                                        		<option value="Aragua"
		                                        			class="hide c16"
		                                        			>Aragua</option>
		                                        	
		                                        		<option value="Apure"
		                                        			class="hide c16"
		                                        			>Apure</option>
		                                        	
		                                        		<option value="Carabobo"
		                                        			class="hide c16"
		                                        			>Carabobo</option>
		                                        	
		                                        		<option value="Caracas"
		                                        			class="hide c16"
		                                        			>Caracas</option>
		                                        	
		                                        		<option value="Bolivar"
		                                        			class="hide c16"
		                                        			>Bolivar</option>
		                                        	
		                                        		<option value="Falcon"
		                                        			class="hide c16"
		                                        			>Falcon</option>
		                                        	
		                                        		<option value="Lara"
		                                        			class="hide c16"
		                                        			>Lara</option>
		                                        	
		                                        		<option value="Marida"
		                                        			class="hide c16"
		                                        			>Marida</option>
		                                        	
		                                        		<option value="Sucre"
		                                        			class="hide c16"
		                                        			>Sucre</option>
		                                        	
		                                        		<option value="Tachira"
		                                        			class="hide c16"
		                                        			>Tachira</option>
		                                        	
		                                        		<option value="Zulia"
		                                        			class="hide c16"
		                                        			>Zulia</option>
		                                        	
	                                        	
											</select>
										</div>
										<a href="/ciudades" class="moreLink">Ver más ciudades</a>
									</div>
								</div>
								<button class="btn-action blueBtn">Listo</button>
							</form>
						</div>
					</div>
				</li>

				
			</ul>
		</div>
	</div>
</header>



		<!--Home background-->
		<section class="homeBg">
			<div class="parallaxImageContainer">
				<img src="http://placehold.it/1932×1280" data-index="0"
					style="transform: translate3d(0px, -447px, 0px); opacity: 1;">
			</div>
			<div class="home-gradient"></div>
			<!--categorias top-->
			



<ul class="TopCategories">
	<li>
		
		<a href="http://www.paginasamarillas.com.sv/servicios/moteles" rel="Index,Follow" title="Moteles">
			<span class="icon-pa_49"></span>&nbsp;Moteles
		</a>
	</li>
	<li>
		
		<a href="http://www.paginasamarillas.com.sv/servicios/cooperativas" rel="Index,Follow" title="Cooperativas">
			<span class="icon-pa_52"></span>&nbsp;Cooperativas
		</a>
	</li>
	<li>
		
		<a href="http://www.paginasamarillas.com.sv/servicios/restaurantes" rel="Index,Follow" title="Restaurantes">
			<span class="icon-pa_07"></span>&nbsp;Restaurantes
		</a>
	</li>
	<li>
		
		<a href="http://www.paginasamarillas.com.sv/servicios/mariachis" rel="Index,Follow" title="Mariachis">
			<span class="icon-pa_53"></span>&nbsp;Mariachis
		</a>
    </li>
	<li>
		
		<a href="http://www.paginasamarillas.com.sv/servicios/taxis" rel="Index,Follow" title="Taxis">
			<span class="icon-pa_58"></span>&nbsp;Taxis
		</a>
	</li>
</ul>
		</section>
				
		
		
		
		
			<section >
				<!--modulo de conversión-->

				
		</section>
		

		

    </section>

		


	<!--Modulo contenido-->
	<section id="seccion_articulos">
		<div class="container contentWrap">

			<div class="title">
				Artículos <b>recomendados</b>
			</div>
			
		<div class="row contentPost">
         
         		<div class="col-md-2">
         				<div class="contentDate">
							<span class="cat-1 semibold cat-a">Automotriz</span>  
						</div>
								
						<div class="contentImg">
							<a href="/automotriz/todas" rel="nofollow"> 
								<img src="/view/global/common/images/content/IMG-Automotriz-01.jpg" alt="Automotriz" title="">
							</a>
						</div>
						<div class="contentBox">
							<div>								
								<div class="description" data-description="">
									Noticias, eventos, consejos de mantenimiento y los m&acute;s recientes avances tecnol&oacute;gicos en la industria automotriz.
								</div>
								<a href="/automotriz/todas" class="moreLink" rel="nofollow">
									Ver contenidos
								</a>
							</div>
						</div>
					</div>
					<div class="col-md-2">
						<div class="contentDate">
							<span class="cat-1 semibold cat-ed">Educaci&oacute;n</span>  
						</div>
								
						<div class="contentImg">
							<a href="/educacion/todas" rel="nofollow"> 
								<img src="/view/global/common/images/content/IMG-Educacion-01.jpg" alt="Educacion" title="">
							</a>
						</div>
						<div class="contentBox">
							<div>
								<div class="description" data-description="">
									Cursos, becas, t&eacute;cnicas de estudio, informaci&oacute;n laboral y todos los avances del sector educativo.
								</div>
								<a href="/educacion/todas" class="moreLink" rel="nofollow">
									Ver contenidos
								</a>
							</div>
						</div>
					</div>
				
					<div class="col-md-2">
						<div class="contentDate">
							<span class="cat-1 semibold cat-ch">Casa y hogar</span>  
						</div>
						<div class="contentImg">
							<a href="/casa-y-hogar/todas" rel="nofollow"> 
								<img src="/view/global/common/images/content/IMG-Hogar-01.jpg" alt="Casa y Hogar" title="">
							</a>
						</div>
						<div class="contentBox">
							<div>
								<div class="description" data-description="">
									Tendencias innovadoras, recetas de cocina y &uacute;tiles pr&aacute;cticas para el  bienestar del hogar.
								</div>
								<a href="/casa-y-hogar/todas" class="moreLink" rel="nofollow">
									Ver contenidos
								</a>
							</div>
						</div>
					</div>
				
					<div class="col-md-2">
						<div class="contentDate">
							<span class="cat-1 semibold cat-m">Mascotas</span>  
						</div>
								
						<div class="contentImg">
							<a href="/mascotas/todas" rel="nofollow"> 
								<img src="/view/global/common/images/content/IMG-Mascotas-01.jpg" alt="Mascotas" title="">
							</a>
						</div>
						<div class="contentBox">
							<div>
								<div class="description" data-description="">
									Consejos de salud, educaci&oacute;n, tips de alimentaci&oacute;n y cuidados para mejorar la calidad de vida de tus mascotas.
								</div>
								<a href="/mascotas/todas" class="moreLink" rel="nofollow" >
									Ver contenidos
								</a>
							</div>
						</div>
					</div>
				
					<div class="col-md-2">
						<div class="contentDate">
								<span class="cat-1 semibold cat-m">Estilo de vida</span>  
						</div>
								
						<div class="contentImg">
							<a href="/estilo-de-vida/todas" rel="nofollow"> 
								<img src="/view/global/common/images/content/IMG-Estilo-01.jpg" alt="Estilo de vida" title="">
							</a>
						</div>
						<div class="contentBox">
							<div>
							
								<div class="description" data-description="">
									Destinos tur&iacute;sticos, opciones gastron&oacute;micas, actividades de entretenimiento y consejos para una llevar una vida saludable.
								</div>
								<a href="/estilo-de-vida/todas" class="moreLink" rel="nofollow" >
									Ver contenidos
								</a>
							</div>
						</div>
					</div>
				
					
				

			</div>
		</div>
	</section>


		<!--Modulo App-->
		<section class="descarga-app">
			
			<a href="/movil" target="_blank" class="link_app"></a>			
				<div class="container">
					<div class="col-md-8 col-lg-8 padding-off">
						<div class="title">
							Descarga nuestro <b>aplicativo móvil</b>
						</div>
						<p class="subtitle">
							Con la App de Páginas Amarillas encuentra información precisa de los establecimientos comerciales más cercanos a tu ubicación. Descárgala desde Play Store o App Store.
						</p>
						<div class="app-buttons">
							<a target="_blank" href="https://play.google.com/store/apps/details?id=com.paginasamarillas&feature=search_result"
								class="btn pa-icon icon-googleplay"></a> <a target="_blank"
								href="https://itunes.apple.com/co/app/paginas-amarillas/id455440191?mt=8" class="btn pa-icon icon-appstore"></a>
						</div>
						<div class="gradientSocial"></div>
					</div>
				</div>
			
		</section>
	

		<!-- TODO QUEMADO para salida de Ecuador -->

	<!-- 	
		 
		<!-- TODO QUEMADO para salida de Guatemala -->
		
		 
				


<!-- secciones más buscadas-->
<section>


	<div class="container sectionWrap">

        <h2 class="title">
            Secciones <b>más buscadas</b>
         </h2>

	 <ul class="listWrap row">
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/clubes-nocturnos">Clubes nocturnos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/ferreterias">Ferreter&iacute;as en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/colegios">Colegios en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/floristerias">Florister&iacute;as en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/hoteles">Hoteles en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/abogados">Abogados en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/bancos">Bancos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/laboratorios-clinicos">Laboratorios cl&iacute;nicos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/farmacias">Farmacias en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/salones-de-belleza">Salones de belleza en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/repuestos-para-vehiculos">Repuestos para veh&iacute;culos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/maquila">Maquila en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/armas-de-fuego">Armas de fuego en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/cerrajerias">Cerrajer&iacute;as en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/librerias">Librer&iacute;as en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/clinicas-veterinarias">Cl&iacute;nicas veterinarias en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/imprentas">Imprentas en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/laboratorios-farmaceuticos">Laboratorios farmac&eacute;uticos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/ginecologia">Ginecolog&iacute;a en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/dentistas">Dentistas en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/telefonos">Tel&eacute;fonos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/reciclaje">Reciclaje en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/panaderias">Panader&iacute;as en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/agencias-de-viajes">Agencias de viajes en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/talleres-de-mecanica-automotriz">Talleres de mec&aacute;nica automotriz en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/clinicas">Cl&iacute;nicas en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/alquiler-de-automotores">Alquiler de automotores en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/escuelas-de-idiomas">Escuelas de idiomas en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/productos-lacteos">Productos l&aacute;cteos en San salvador</a>
           		</li>
           	
           	
           		
             	
           		
           		<li class="">
           			
           			
           			
           		
           			<a href="/san-salvador/servicios/gruas">Gr&uacute;as en San salvador</a>
           		</li>
           	
		</ul> 
	</div>

</section>

				
	<!-- Chat servicio al cliente -->
	
			<!-- BEGIN ProvideSupport.com Graphics Chat Button Code -->
			<div id="ci4s1g" class="chatci"></div>
			<div id="sc4s1g" class="chatlive"></div>
			<div id="sd4s1g" class="is-totally-hidden"></div>
			
			<script type="text/javascript">
				var se4s1g=document.createElement("script");
				se4s1g.type="text/javascript";
				var se4s1gs=(location.protocol.indexOf("https")==0?"https":"http")+"://image.providesupport.com/js/0j6pz2c2mgcat1957t79e76sti/safe-standard.js?ps_h=4s1g&ps_t="+new Date().getTime();
				setTimeout("se4s1g.src=se4s1gs;document.getElementById('sd4s1g').appendChild(se4s1g)",1)
			</script>
			<noscript><div style="display:inline"><a href="http://www.providesupport.com?messenger=0j6pz2c2mgcat1957t79e76sti">Live Chat</a></div></noscript>
			<!-- END ProvideSupport.com Graphics Chat Button Code -->
		
	

	<!-- Footer -->
	

<footer>
    <!--footer tags-->
    <div class="tagWrap row margin-off">
        <ul class="col-lg-12 col-md-12 col-sm-12 menu-tags">
            <li>
                <a href="http://publitag.co" target="_blank"><i class="icon-pa_12"></i>Publitags</a>
            </li>
            <li>
                <a href="https://www.publicar.com/servicio-al-cliente/preguntas-frecuentes-cuentas-correo" target="_blank"><i class="icon-pa_13"></i>Webmail</a>
            </li>
            <li>
                <a href="/movil" target="_blank"><i class="icon-pa_14"></i>App</a>
            </li>
            <li>
                <a onclick="return clickGuidePrinted(this,TipoClick.CLIC_WEB,Pagina.PAGE_HOME);" href="http://sites.paginasamarillas.com/directorio/home.html" target="_blank"><i class="icon-pa_16"></i>Directorios</a>
            </li>
            <li>
                <span class="is-link" data-toggle="modal" data-target="#anuncia-modal"><i class="icon-pa_15"></i>Anúnciate</span>
            </li>
            <li>
                <span class="is-link" data-toggle="modal" data-target="#updateInfoModal"><i class="icon-pa_17"></i>Actualizar información</span>
            </li>
            <li>
                <a href="http://www.publicar.com/unidadessac" target="_blank"><i class="icon-pa_18"></i>Servicio al Cliente</a>
            </li>
            <li>
                <a href="/mapa-del-sitio"><i class="icon-pa_19"></i>Mapa del Sitio</a>
            </li>
            <li>
                <a href="/ayuda"><i class="icon-pa_73"></i>Ayuda</a>
            </li>
        </ul>
    </div>
    <div class="seoWrap container">
        <div class="row">
            <div class="col-md-5">
                <div class="titleFooter">Otros de nuestros sitios</div>
                <ul class="sitesList">
                    <li><a href="http://www.publicar.com/" target="_blank">Publicar</a></li>
                    <li><a href="http://www.publicar.com/blog/" target="_blank">Visite nuestro blog</a></li>
                    <li><a href="http://www.publicar.com/marketing-directo?hs_preview=xkh0kjfn-1911279459" target="_blank">Contacto inteligente</a></li>
                    <li><a href="http://www.ciudadguru.com.sv/" target="_blank">Ciudad Gurú</a></li>
                    <li><a href="http://www.gurucasayhogar.com.sv/" target="_blank">Gurú Casa y Hogar</a></li>
                    <li><a href="http://www.guruautomotriz.com.sv/" target="_blank">Gurú Automotriz</a></li>
					<li><a href="http://www.gurumascotas.com.sv/" target="_blank">Gurú Mascotas</a></li>
                    <li><a href="http://www.gurueducacion.com.sv/" target="_blank">Gurú Educación</a></li>
                    <li><a href="http://www.gurukids.com.sv/" target="_blank">Gurú Kids</a></li>
                    <li><a href="http://www.gurusalud.com.sv/" target="_blank">Gurú Salud</a></li>
                </ul>
            </div>
            <div class="col-md-5">
                <div class="titleFooter">Contenido</div>
               
                <p class="contentTxt ctxt">
                P&aacute;ginas Amarillas es el directorio m&aacute;s grande de Latinoam&eacute;rica, en el que encontrar&aacute;s la solución que necesitas de forma r&aacute;pida y sencilla. Realiza tus b&uacute;squedas comerciales desde cualquier lugar y dispositivo.
                </p>
            </div>
            <div class="col-md-2">
                <div class="titleFooter">S&iacute;guenos</div>
                <ul class="footNetwork">
                    <li><a href="https://www.facebook.com/PaginasAmarillasSV" target="_blank"><i class="pa-icon icon-fb"></i></a></li>
                    <li><a href="https://twitter.com/PublicarCol" target="_blank"><i class="pa-icon icon-tw"></i></a></li>
                    <li><a href="https://www.youtube.com/user/PaginasAmarillasSV" target="_blank"><i class="pa-icon icon-yt"></i></a></li>
                </ul>
                <span class="is-link moreLink" onclick="guru.commons.setDesktopCookie()">
                    Versión móvil <span class="icon-pa_01"></span>
                </span>
            </div>
        </div>
        <div class="row">
            <div class="col-md-8 pull-left">
                <div class="titleFooter">Protección de datos personales</div>
                <p class="contentTxt">
                    La política de tratamiento de datos personales de Publicar puede ser consultada&nbsp;<a href="https://www.publicar.com/manejo-datos" target="_blank">aquí.</a>
                </p>
            </div>
        </div>
         <hr>
        <div class="row legales">
            <div class="col-md-12">
                <p>El portal de negocios de PaginasAmarillas.com de Publicar contiene la información comercial de 15 países de Latinoamérica.</p>
                <p>
                	Todas las marcas registradas son propiedad de la compañía respectiva o de Publicar. La reproducción total o parcial de cualquier material contenido en este portal está prohibido.&nbsp;<a href="/aviso-legal">AVISO LEGAL</a>&nbsp;©Copyright&nbsp;2018
                </p>
                <br>
               
            </div>
        </div>
    </div>
</footer>
	


<div id="scrolltop" class="icon-pa_42"></div>

<script>
	var COUNTRY = "sv",
		COUNTRY_NAME = "El Salvador",
		GLOBAL_HOME_PATH = "http://www.paginasamarillas.com.sv",
		GLOBAL_SUB_DOMAIN = "www.paginasamarillas.com.sv",
		GLOBAL_KEYWORD = "",
		GLOBAL_LOCALITY = "",
		GLOBAL_SEARCHTYPE = "",
		GLOBAL_MOBILE_PATH = "http://m.paginasamarillas.com.sv",
		CITY = "",
		RECAPTCHA_ID = '6Ldi1CgTAAAAACT6EyFR8xxSN_FyFcj0omehH2QZ';
		//para yell-analytics
		FORBIDDEN_WORDS = 'erotica;sex;scorts;masajes;masaje;prepago;prepagos;acompañante;acompanante;acompañantes;acompanantes;masajistas;masajista;articulos para adultos;artículos para adultos;articulos eroticos;artículos eróticos;eróticos;erotico;eroticos;abusador;abusadora;abuso;abusos;adulterio;agujero;agujeros;anal;anales;androgeno;androgenos;ano;bálano;bestialidad;Bisexual;bisexuales;bondage;bubbie;bubbies;busto;bustos;cachondear;cachondo;caliente;carnal;carnales;chocho;chupada;chupadas;chupar;Cita;Citas;clitoris;coito;Colegiala;colegialas;condon;condones;conejita;conejito;consolador;consoladores;coño;coños;copula;copular;cornuda;cornudas;cornudo;cornudos;culo;culos;desnudismo;desnudos;duro;erótica;erótico;erotismo;esperma;espermas;extasis;eyaculación;eyaculaciones;eyacular;falo;falos;fetichismo;follar;fornicador;fornicadores;fornicar;Gay;gemido;gemidos;genitales;gigolo;gigolos;glande;glandes;Hermafrodita;hermafroditas;himen;Homosexual;homosexuales;incesto;joder;lame;lamer;lascivo;lascivos;lechita;lechoso;lechosos;lesbia;Lesbiana;lesbianas;libido;lujuria;lujurias;lujuriosa;lujuriosas;lujurioso;lujuriosos;maduro;mamada;mamadas;mamar;maricón;Masturbación;Menores;mierda;mierdas;Motel;Moteles;mujerzuela;mujerzuelas;munequita;muñeca;muñecas;Necrofilia;negra;negro;obsceno;obsenidades;orgía;orgías;pecho;pechos;Pedofilia;pene;penes;perra;pezón;pezones;pipi;pipis;polla;porno;pornografia;prepucio;prepucios;preservativo;preservativos;promiscuo;promiscuos;prostituta;prostitutas;pulpa;puta;putas;puto;putos;ramera;rameras;sádico;sádicos;sadomasoquismo;sadomasoquista;sadomasoquistas;sapo;seducción;seducciones;seducir;semen;seminal;sensual;sensuales;sexo;sexual;sexuales;sexualidad;sexy;snuff;swinger;tetas;Trío;vagina;vaginas;verga;vergas;vibradores;violación;violaciones;violador;violadora;virgen;virgenes;virgo;viril;voyerismo;voyeur;vulva;zorra;hidromasajes;masajes terapeuticos;masaje terapeutico;ofisex;unisex;sexta;sexto;sextinvalle;sexteto;sextiri;sexiquartz;isex;asexma;sexco;disexport;gasexpress;juegosextremos.com;misex;sexi jeans;gasex';
		guru = [];

	//textos internacionalizados para el suggest
	var suggestText = {
			titleWhatLeft: 	'Secciones',
			titleWhatRight: 'Empresas',
			titleWhereLeft:	'Ciudades',
			titleWhereRight:'Estado',
			errorWhatLeft:	'No se han encontrado secciones',
			errorWhatRight:	'No se han encontrado empresas',
	};
</script>



	<script>var TIMEZONE = -6;</script>




<!-- jQuery (necessary for Bootstrap's JavaScript plugins) -->
<!--<script src="https://ajax.googleapis.com/ajax/libs/jquery/1.12.4/jquery.min.js"></script> -->

<!-- Modulo Actualizar Datos -->


<div id="updateInfoModal" class="modal fade modal-guru" tabindex="-1"
	role="dialog" aria-labelledby="myLargeModalLabel">
	<div class="modal-dialog" role="document">
		<div class="modal-content">
			<div class="modal-header">
				<button type="button" class="close" data-dismiss="modal" aria-label="Close">
					<span aria-hidden="true">×</span>
				</button>
			</div>
			<div class="modal-body background-actualizainfo" data-mod-body data-steps-container>
				<form id="updateInfoForm" action="/sendMailInfoUpdate.action" data-mod-form novalidate>
					<input type="hidden" name="country" value="El Salvador">
					<input type="hidden" name="mailtype" value="3">

					<div>
						<!--titulo-->
						<div class="title">
							<span class="titleBold">Actualiza tu información</span>
						</div>
						<p>Los campos marcados con * son obligatorios</p>
					</div>
					
					<div class="row contactFormWrap">
						<div class="col-xs-12 bold">
							Información personal
						</div>

						<div class="col-xs-12 col-sm-5 required">
							<label for="actualizaFullName">Nombres y Apellidos</label>
							<input id="actualizaFullName" name="FullName" type="text" placeholder="Ingresa tu nombre completo" required>
							<div class="error hide">Su Nombre es obligatorio</div>
						</div>
						<div class="col-xs-12 col-sm-5 required">
							<label for="actualizaupdatephone">Número de contacto</label>
							<input id="actualizaupdatephone" name="updatephone" type="number" placeholder="Ej. 312 555 2342" required>
							<div class="error hide">Su Número de contacto es obligatorio</div>
						</div>
						<div class="col-xs-12 col-sm-5 required">
							<label for="actualizaid">Tipo y Número de documento</label>
							<div class="row">
								<div class="col-xs-4 padding-right-off selectWrap">
									<select name="typeId" class="anunciaSelect">
										<option value="CC">CC</option>
										<option value="CE">CE</option>
										<option value="DI">DI</option>
									</select>
								</div>
								<div class="col-xs-8 required">
									<input id="actualizaid" name="id" type="number" placeholder="Ej:1020764824" required>
									<div class="error hide">Su número y tipo de identificación son obligatorios.</div>
								</div>
							</div>
						</div>
						<div class="col-xs-12 col-sm-5 required">
							<label for="actualizaCity">Ciudad</label>
							<input id="actualizaCity" name="City" type="text" placeholder="Ej.San Juan" required  data-suggest="location" autocomplete="off">
							<div class="error hide">Ingrese la ciudad</div>
							<div id="actualizaCityList" class="sections-list hide"></div>
						</div>
						<div class="col-xs-12 col-sm-10 required">
							<label for="actualizaCompanyName">Nombre de tu empresa</label>
							<input id="actualizaCompanyName" name="CompanyName" type="text" placeholder="Ej.Hotel Sauces" required>
							<div class="error hide">El nombre de la empresa es obligatorio.</div>
						</div>
						
						<div class="col-xs-12 col-sm-10 required">
							<label for="actualizaemail">Email</label>
							<input id="actualizaemail" name="email" type="email" placeholder="Ej.nombreusuario@emmail.com" required>
							<div class="error hide">Su correo electrónico es obligatorio.</div>
						</div>
						<div class="col-xs-12 col-sm-10">
							<label for="actualizacomment">Dejanos tu comentario</label> 
							<textarea id="actualizacomment" name="Comments" placeholder="Escribe tu inquietud a Pizza Piccolo" maxlength="1024"  aria-invalid="true"></textarea>
						</div>

						<div class=" col-xs-12 col-sm-10 form-legal required">
        					<input name="terms" type="checkbox" required>
		        			<p>Conozco y acepto&nbsp;<a target="_blank" href="/aviso-legal">términos y condiciones</a>&nbsp; y el tratamiento de mis datos personales de conformidad con la Política de&nbsp; 
		        			<a target="_blank" href="https://www.publicar.com/manejo-datos">Tratamiento de Datos Personales</a>&nbsp;y el&nbsp; <a target="_blank" href="https://www.publicar.com/manejo-datos" >&nbsp;Aviso de Privacidad&nbsp;</a>&nbsp;de Publicar.</p>
        					<div class="error hide">Debe aceptar los términos y condiciones.</div>
       					</div>
						<div class="col-xs-12 col-sm-10">
							<div id="updateInfoError"></div>
						</div>
						<div class="col-xs-12 col-sm-10">
							<button class="btn-more contactLite pull-left">Enviar</button>
						</div>
							
					</div>
				</form>

				<div class="result-message hide">
					<div class="message-ok">
						<div class="title">Gracias por actualizar <b class="titleBold">tus datos. </b></div>
						<p>Pronto nos pondremos en contacto contigo para verificar que estos <b>sean correctos.</b></p>
					</div>
					<div class="message-error">
						<div class="title">Se ha producido un <b>error</b></div>
						<p>Por favor, espere un momento e intente nuevamente</p>
					</div>
					<div class="btn-action blueBtn" data-dismiss="modal" aria-label="Close" data-mod-reset>Listo</div>
				</div>
			</div>
		</div>
	</div>
</div>



<!-- Modulo confirmar edad -->


<div id="edadModal" class="modal fade modal-guru" tabindex="-1"
	role="dialog" aria-labelledby="myLargeModalLabel">
	<div class="modal-dialog" role="document">
		<div class="modal-content">
			<div class="modal-header">
				<button type="button" class="close" data-dismiss="modal" aria-label="Close">
					<span aria-hidden="true">×</span>
				</button>
			</div>
			<div class="modal-body background-edad" data-mod-body data-steps-container>
				<div class="result-message">
					<div>
						<div class="title">Confírmanos <b>tu edad.</b></div>
						<p>Manifiesto ser mayor de edad y que ingreso a este sitio web y a su contenido <b>bajo mi esclusiva responsabilidad</b>.Soy consciente de que en este sitio es posible encontrar contenidos de naturaleza sexual al cual accedo de manera voluntaria.</p>
					</div>
					<div>
						<div id="age_invalid" class="btn btn-action greyBtn ">Soy menor de 18 años</div>
						<div id="age_valid" class="btn btn-action blueBtn">Soy mayor de 18 años</div>
					</div>
				</div>
			</div>
		</div>
	</div>
</div>



<!-- Anuncia -->

<div id="anuncia-modal" class="modal fade modal-guru" tabindex="-1"
	role="dialog" aria-labelledby="myLargeModalLabel">
	<div class="modal-dialog " role="document">
		<div class="modal-content">
			<div class="modal-header">
				<button type="button" class="close" data-dismiss="modal"
					aria-label="Close">
					<span aria-hidden="true">×</span>
				</button>
			</div>
			<div class="modal-body background-anuncia anuncia-hbspt" data-mod-body data-steps-container>
				
				
					<div class="title">
						<b>Anúnciate</b>
					</div>
					<p class="text-title">
						Los campos marcados con * son obligatorios
					</p>
			
					<script charset="utf-8" type="text/javascript" src="//js.hsforms.net/forms/v2.js"></script>
					
					<script>
						hbspt.forms.create({
							sfdcCampaignId: '701f1000001cKyCAAU',
							portalId: '251261',
							formId: '3eb6590b-dcd4-413e-b46e-d7ab6b0cefa0'
						});
					</script>

					<style>
						#anuncia-modal .message-ok{
						display:block;
						}
						.submitted-message{
							color: #000;
						    font-size: 33px;
						    line-height: 32px;
						    margin-bottom: 10px;
						    margin-top: 30px;
						   	font-family: 'SourceSansProRegular';
						}
						
					</style>
					<div class="message-ok">
						<p>
							Gracias por hacer parte del directorio electrónico más completo y confiable de América Latina. </br> Pronto nos pondremos en contacto contigo para finalizar el proceso de inscripción.
						</p>   
                      <br />
                      
                      <div class="btn-action btn-ready blueBtn" >Listo</div>
                      </div>

                    
					<script>
					$('#anuncia-modal .message-ok').hide();
					var checkExist = setInterval(function() {
						if ($(".submitted-message").length > 0) {
							$('#anuncia-modal .title').hide();
							$('#anuncia-modal .text-title').hide();
							$('#anuncia-modal .message-ok').show();
						}
						}, 100); // check every 100ms
					
					$('#anuncia-modal .btn-ready').click(function() {
					    location.reload();
					});
					</script>
				
			</div>
		</div>
	</div>
</div>
<script>
/* $(document).bind('DOMNodeInserted', function(e) {
	
		$( ".submitted-message" ).html( "<div class='message-ok'> <div class='title'>Gracias por actualizar <b class='titleBold'>tus datos. </b></div><p>Pronto nos pondremos en contacto contigo para verificar que estos <b>sean correctos.</b></p></div><div class='btn-action blueBtn' data-dismiss='modal' aria-label='Close' data-mod-reset=''>Listo</div>" );
		console.log('cambios dom');
}); */
</script>

<!-- Include all compiled plugins (below), or include individual files as needed -->
<script src="/view/global/common/vendor/bootstrap/js/bootstrap.min.js"></script>
<script src="/view/global/common/vendor/jquery/jquery.cookie.min.js"></script>
<script src="/view/global/common/vendor/js.cookie.js"></script>
<script src="/view/global/common/js/cookies_utils.js"></script>
<script src="/view/global/common/js/modulosCommons.js?20171026"></script>
<script src="/view/global/common/js/commons.js?20171117"></script>
<script src="/view/global/common/js/suggest.js?20170919"></script>
<script src="/view/global/common/js/submit.js?20170831"></script>

<!-- SSO -->

	<script src="/view/global/common/js/index.js?20170906"></script>
	<script src="/view/global/common/js/quotations.js"></script>

	
    



    
   

</body>

</html>