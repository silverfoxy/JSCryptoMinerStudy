


 


 <!DOCTYPE html>
<html lang="en">
    <head>
        <meta charset="utf-8">
        <meta http-equiv="X-UA-Compatible" content="IE=edge">
        <meta name="viewport" content="width=device-width, initial-scale=1">
        <title>Universidad Centroamericana José Simeón Cañas</title>
        <meta name="description" lang="es" content="Universidad para el cambio social, educación superior, calidad educativa, universidad jesuita">
        <meta name="keywords" lang="es" content="Educación, Universidad, Pregrados, Postgrados, Desarrollo estudiantil, vida universitaria, mártires, cursos libres, admisión, uca, El Salvador, martires uca,Investigación, investigadores, investigaciones, responsabilidad social universitaria, responsabilidad social, ausjal, teologia de la liberacion, teología de la liberación, jon sobrino, Ignacio Ellacuría" />
        <meta name="author" content="UCA - www.uca.edu.sv" />
        <meta name="robots" content="index,follow" />
        <meta name="revisit-after" content="1 days" />
        <meta http-equiv="Cache-Control" content="no-cache"> 
        <meta http-equiv="Expires" content="0"> 
        <meta http-equiv="Pragma" content="no-cache">
        <link href="http://www.uca.edu.sv/wp-content/themes/kubo/css/bootstrap.min.3.2.0.css?15438051" rel="stylesheet"> 
        <link href="http://www.uca.edu.sv/wp-content/themes/kubo/css/tema.css?487518371" rel="stylesheet">
        <link href="http://www.uca.edu.sv/wp-content/themes/kubo/css/bootstrap-responsive-tabs.css" rel="stylesheet">   
        <!--[if lt IE 9]>
          <script src="https://oss.maxcdn.com/html5shiv/3.7.3/html5shiv.min.js"></script>
          <script src="https://oss.maxcdn.com/respond/1.4.2/respond.min.js"></script>
        <![endif]-->
        <script src='https://www.google.com/recaptcha/api.js'></script>
        <meta name='robots' content='noindex,follow' />
<link rel='dns-prefetch' href='//s.w.org' />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/www.uca.edu.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.7.3"}};
			!function(a,b,c){function d(a){var b,c,d,e,f=String.fromCharCode;if(!k||!k.fillText)return!1;switch(k.clearRect(0,0,j.width,j.height),k.textBaseline="top",k.font="600 32px Arial",a){case"flag":return k.fillText(f(55356,56826,55356,56819),0,0),!(j.toDataURL().length<3e3)&&(k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,65039,8205,55356,57096),0,0),b=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,55356,57096),0,0),c=j.toDataURL(),b!==c);case"emoji4":return k.fillText(f(55357,56425,55356,57341,8205,55357,56507),0,0),d=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55357,56425,55356,57341,55357,56507),0,0),e=j.toDataURL(),d!==e}return!1}function e(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var f,g,h,i,j=b.createElement("canvas"),k=j.getContext&&j.getContext("2d");for(i=Array("flag","emoji4"),c.supports={everything:!0,everythingExceptFlag:!0},h=0;h<i.length;h++)c.supports[i[h]]=d(i[h]),c.supports.everything=c.supports.everything&&c.supports[i[h]],"flag"!==i[h]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[i[h]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(g=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",g,!1),a.addEventListener("load",g,!1)):(a.attachEvent("onload",g),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),f=c.source||{},f.concatemoji?e(f.concatemoji):f.wpemoji&&f.twemoji&&(e(f.twemoji),e(f.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='https://api.w.org/' href='http://www.uca.edu.sv/wp-json/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://www.uca.edu.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://www.uca.edu.sv/wp-includes/wlwmanifest.xml" /> 
<meta name="generator" content="WordPress 4.7.3" />
        <script type="text/javascript">

        var _gaq = _gaq || [];
        _gaq.push(['_setAccount', 'UA-27456897-1']);
        _gaq.push(['_trackPageview']);

        (function() {
        var ga = document.createElement('script'); ga.type = 'text/javascript'; ga.async = true;
        ga.src = ('https:' == document.location.protocol ? 'https://ssl' : 'http://www') + '.google-analytics.com/ga.js';
        var s = document.getElementsByTagName('script')[0]; s.parentNode.insertBefore(ga, s);
        })();

        </script>
    </head>
<body id="main">
    <div id="mySidenav" class="sidenav">
        <a href="javascript:void(0)" class="closebtn" onclick="closeNav()">&times;</a>
        <a href="http://www.uca.edu.sv/noticias/">Noticias UCA</a>
        <a href="http://abaco.uca.edu.sv/bfi/">Biblioteca P. Idoate</a>
        <a href="http://bibteol.uca.edu.sv/">Biblioteca de Teología</a>
        <a href="http://www.uca.edu.sv/cartelera/">Cartelera</a>
        <a href="http://www.uca.edu.sv/calendario-academico/">Calendario académico</a>       
        <a href="http://www.uca.edu.sv/personal/" target="_ventana">Directorio</a>             
    </div>
    <header>
        <div class="menu-layer hidden-xs">
        <div class="container-fluid no-padding fondo-1 hidden-xs">
            <button type="button" class="menuGeneralUCA" id="menuGeneralUCA" >
            <span class="icon-bar-UCA"></span>
            <span class="icon-bar-UCA"></span>
            <span class="icon-bar-UCA"></span>
        </button><div class="menuGeneral"><ul id="menu-menu-lateral" class="MenuG"><li id="menu-item-3796" class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home current-menu-ancestor current-menu-parent menu-item-has-children menu-item-3796 dropdown active"><a title="Inicio" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Inicio <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-3797" class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-3797 active"><a title="Eventos y noticias" href="http://www.uca.edu.sv/#eventos-noticias">Eventos y noticias</a></li>
	<li id="menu-item-3798" class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-3798 active"><a title="Lo más reciente" href="http://www.uca.edu.sv/#lo-mas-reciente">Lo más reciente</a></li>
	<li id="menu-item-3799" class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-3799 active"><a title="#OrgulloUCA" href="http://www.uca.edu.sv/#orgullo-uca">#OrgulloUCA</a></li>
</ul>
</li>
<li id="menu-item-3800" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children menu-item-3800 dropdown"><a title="Nuevo ingreso y admisión" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Nuevo ingreso y admisión <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-3802" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3802"><a title="Pasos" href="http://www.uca.edu.sv/pasos-para-nuevo-ingreso/">Pasos</a></li>
	<li id="menu-item-3803" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3803"><a title="Inscripción a pruebas" href="http://www.uca.edu.sv/admisiones/#inscripcion-pruebas-admision-ciclo-02-2018">Inscripción a pruebas</a></li>
	<li id="menu-item-3804" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3804"><a title="Becas, cuotas y formas de ingreso" href="http://www.uca.edu.sv/admisiones/#becas-cuotas-y-formas-de-ingreso">Becas, cuotas y formas de ingreso</a></li>
	<li id="menu-item-4235" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-4235"><a title="Oferta académica Ciclo 02/2018" href="http://www.uca.edu.sv/admisiones/#oferta-academica-ciclo-02-2018">Oferta académica Ciclo 02/2018</a></li>
	<li id="menu-item-3805" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3805"><a title="Carreras y diagnóstico vocacional" href="http://www.uca.edu.sv/admisiones/#conoce-nuestras-carreras-y-encuentra-tu-vocacion">Carreras y diagnóstico vocacional</a></li>
	<li id="menu-item-3806" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3806"><a title="¿Necesitas más ayuda?" href="http://www.uca.edu.sv/admisiones/#necesitas-mas-ayuda">¿Necesitas más ayuda?</a></li>
</ul>
</li>
<li id="menu-item-3809" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children menu-item-3809 dropdown"><a title="Oferta académica" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Oferta académica <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-3814" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3814"><a title="Carreras" href="http://www.uca.edu.sv/oferta-academica/carreras/">Carreras</a></li>
	<li id="menu-item-3815" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3815"><a title="Maestrías y doctorados" href="http://www.uca.edu.sv/postgrados/">Maestrías y doctorados</a></li>
	<li id="menu-item-3816" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3816"><a title="Formación continua" href="http://www.uca.edu.sv/formacion-continua/">Formación continua</a></li>
	<li id="menu-item-3817" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3817"><a title="Cursos de idiomas" href="http://www.uca.edu.sv/escuela-de-idiomas/">Cursos de idiomas</a></li>
</ul>
</li>
<li id="menu-item-3818" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children menu-item-3818 dropdown"><a title="Vida estudiantil" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Vida estudiantil <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-3940" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3940"><a title="Ciclo 01/2018" href="http://www.uca.edu.sv/vida-estudiantil/#ciclo-01-2018">Ciclo 01/2018</a></li>
	<li id="menu-item-3819" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3819"><a title="Evaluación a docentes Ciclo 03/2017" href="http://www.uca.edu.sv/vida-estudiantil/#evaluacion-en-linea-a-docentes-ciclo-032017">Evaluación a docentes Ciclo 03/2017</a></li>
	<li id="menu-item-3822" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3822"><a title="Ciclo 03/2017 (interciclo)" href="http://www.uca.edu.sv/vida-estudiantil/#ciclo-032017-interciclo">Ciclo 03/2017 (interciclo)</a></li>
	<li id="menu-item-3823" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3823"><a title="Desarrollo estudiantil" href="http://www.uca.edu.sv/vida-estudiantil/#desarrollo-estudiantil">Desarrollo estudiantil</a></li>
</ul>
</li>
<li id="menu-item-4337" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-4337"><a title="Graduados" href="http://www.uca.edu.sv/graduados/">Graduados</a></li>
<li id="menu-item-3824" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3824"><a title="Acerca de la UCA" href="http://www.uca.edu.sv/acerca-de-la-uca/">Acerca de la UCA</a></li>
<li id="menu-item-3825" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3825"><a title="Docencia" href="http://www.uca.edu.sv/acerca-de-la-uca/docencia/">Docencia</a></li>
<li id="menu-item-3826" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3826"><a title="Investigación" href="http://www.uca.edu.sv/acerca-de-la-uca/investigacion/">Investigación</a></li>
<li id="menu-item-3827" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3827"><a title="Proyección social" href="http://www.uca.edu.sv/acerca-de-la-uca/proyeccion-social/">Proyección social</a></li>
<li id="menu-item-3828" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children menu-item-3828 dropdown"><a title="Sobre nosotros" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Sobre nosotros <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-3829" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3829"><a title="Historia" href="http://www.uca.edu.sv/historia/">Historia</a></li>
	<li id="menu-item-3830" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3830"><a title="Misión y visión" href="http://www.uca.edu.sv/mision-y-vision/">Misión y visión</a></li>
	<li id="menu-item-3831" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3831"><a title="Identidad y funciones" href="http://www.uca.edu.sv/identidad-y-funciones/">Identidad y funciones</a></li>
	<li id="menu-item-3832" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3832"><a title="Mártires UCA" href="http://www.uca.edu.sv/biografias-de-los-martires-uca/">Mártires UCA</a></li>
	<li id="menu-item-3833" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3833"><a title="Noticias y editoriales" href="http://www.uca.edu.sv/noticias/">Noticias y editoriales</a></li>
	<li id="menu-item-3834" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3834"><a title="Cartelera informativa" href="http://www.uca.edu.sv/cartelera/">Cartelera informativa</a></li>
	<li id="menu-item-3835" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3835"><a title="Prensa" href="http://www.uca.edu.sv/acerca-de-la-uca/prensa/">Prensa</a></li>
	<li id="menu-item-3836" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3836"><a title="Documentos institucionales" href="http://www.uca.edu.sv/documentos-institucionales/">Documentos institucionales</a></li>
	<li id="menu-item-3837" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3837"><a title="Repositorio Institucional" href="http://repositorio.uca.edu.sv/jspui/">Repositorio Institucional</a></li>
	<li id="menu-item-3838" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3838"><a title="Publicaciones" href="http://www.uca.edu.sv/publicaciones/">Publicaciones</a></li>
</ul>
</li>
<li id="menu-item-3839" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3839"><a title="Servicios" href="http://www.uca.edu.sv/acerca-de-la-uca/#nuestros-servicios">Servicios</a></li>
<li id="menu-item-3840" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-3840"><a title="La UCA en datos" href="http://www.uca.edu.sv/acerca-de-la-uca/#la-uca-en-datos">La UCA en datos</a></li>
</ul></div>            <div class="menu-link padding-top padding-bottom" onclick="openNav()">
                <img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/link-rapidos.png">
            </div>            
            <div class="container">                
                <div class="col-xs-12 col-sm-6 col-md-6  pull-right padding-top padding-bottom text-right">
                    <div class="mail-uca">
                        <a href="http://correo.uca.edu.sv" data-toggle="tooltip" data-placement="bottom" title="Correo institucional">
                            <img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/correo-uca.png" />
                        </a>
                        <a href="https://portal-estudiantes.uca.edu.sv/" data-toggle="tooltip" data-placement="bottom" title="Portal de Estudiantes">
                            <img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/portal-estudiantes.png" />
                        </a>
                        <a href="https://portal-empleados.uca.edu.sv/" data-toggle="tooltip" data-placement="bottom" title="Portal de Empleados">
                            <img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/portal-empleados.png" />
                        </a>


                    </div>
                    <form action="http://www.uca.edu.sv/buscador/" method="get" id="form_bq">
                        <div class="input-group ">
                            <input type="text" class="form-control" placeholder="Buscar" name="q" id="q" value="">
                            <span class="input-group-btn" >
                                <button class="btn btn-default" type="submit"><span class="glyphicon glyphicon-search"></span></button>
                            </span>
                        </div>
                    </form>

       
                </div>
            </div>       
        </div>
        </div>

        <div class="container no-padding barra-movil">
            <nav class="navbar navbar-default  no-margin" role="navigation">
	<div class="navbar-header">
		<button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#menu-uca">
			<span class="sr-only">Toggle navigation</span>
			<span class="icon-bar"></span>
			<span class="icon-bar"></span>
			<span class="icon-bar"></span>
		</button>
		<a class="navbar-brand " href="http://www.uca.edu.sv">
			<div class="logotipo">
				<div class="logo">
					<img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/logo-uca.png" alt="Universidad Centroamericana José Simeón Cañas" title="Universidad Centroamericana José Simeón Cañas" data-toggle="tooltip" data-placement="bottom" class="logo-img">
				</div>
				<div class="logo-texto">
					Universidad Centroamericana<br /> José Simeón Cañas
				</div>
			</div>
		</a>
	    <div class="movil-iconos">
	    	<a href="" data-toggle="modal"  data-target="#comunicaciones">
	    		<!--<span class="glyphicon glyphicon-search fuente-30" data-toggle="tooltip" data-placement="bottom" title="Buscar contenido"></span>-->
	    		<img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/icon-buscar.png" class="img-responsive" style="float:left; margin-right: 5px;" data-toggle="tooltip" data-placement="bottom" title="Buscar contenido" alt="Buscar">
	    	</a> 
	        <a href="http://correo.uca.edu.sv" data-toggle="tooltip" data-placement="bottom" title="Correo institucional">
	            <span class="glyphicon glyphicon-envelope fuente-30" aria-hidden="true"></span>
	        </a>
	    </div>                  
	</div>
	<div id="menu-uca" class="collapse navbar-collapse no-padding"><ul id="menu-menu-1" class="nav navbar-nav navbar-right"><li id="menu-item-600" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-600"><a title="Admisión" href="http://www.uca.edu.sv/admisiones/">Admisión</a></li>
<li id="menu-item-636" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-636"><a title="Oferta académica" href="http://www.uca.edu.sv/oferta-academica/">Oferta académica</a></li>
<li id="menu-item-674" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-674"><a title="Vida estudiantil" href="http://www.uca.edu.sv/vida-estudiantil/">Vida estudiantil</a></li>
<li id="menu-item-683" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-683"><a title="Acerca de la UCA" href="http://www.uca.edu.sv/acerca-de-la-uca/">Acerca de la UCA</a></li>
<li id="menu-item-4336" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-4336"><a title="Graduados" href="http://www.uca.edu.sv/graduados/">Graduados</a></li>
<li id="menu-item-2757" class="hidden-sm hidden-md hidden-lg menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children menu-item-2757 dropdown"><a title="Enlaces directos" href="#" data-toggle="dropdown" class="dropdown-toggle" aria-haspopup="true">Enlaces directos <span class="caret"></span></a>
<ul role="menu" class=" dropdown-menu">
	<li id="menu-item-2771" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2771"><a title="Noticias UCA" href="http://www.uca.edu.sv/noticias/">Noticias UCA</a></li>
	<li id="menu-item-2759" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2759"><a title="Portal de Estudiantes" href="https://portal-estudiantes.uca.edu.sv/">Portal de Estudiantes</a></li>
	<li id="menu-item-2760" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2760"><a title="Portal de Empleados" href="https://portal-empleados.uca.edu.sv/">Portal de Empleados</a></li>
	<li id="menu-item-2756" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2756"><a title="Cartelera" href="http://www.uca.edu.sv/cartelera/">Cartelera</a></li>
	<li id="menu-item-2758" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2758"><a title="Calendario académico" href="http://www.uca.edu.sv/calendario-academico/">Calendario académico</a></li>
	<li id="menu-item-2820" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2820"><a title="Biblioteca P. Idoate" href="http://abaco.uca.edu.sv/bfi/">Biblioteca P. Idoate</a></li>
	<li id="menu-item-2821" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2821"><a title="Biblioteca de Teología" href="http://bibteol.uca.edu.sv/">Biblioteca de Teología</a></li>
	<li id="menu-item-2761" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-2761"><a title="Directorio" href="http://www.uca.edu.sv/personal/">Directorio</a></li>
</ul>
</li>
</ul></div></nav>

        </div>
        <div class="separador"></div>
    </header>
    
    <section>
		
		<div class="container-fluid no-padding">
			<div class="col-md-12 no-padding">
				<div id="banner" class="carousel slide" data-ride="carousel"><div class="carousel-inner anim" role="listbox"><div class='item active'><a href='http://www.uca.edu.sv/admisiones/'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/03/banner-portada-nuevo-ingreso-02-18-3.jpg' alt=''  /></a> 
						<a href='http://www.uca.edu.sv/admisiones/'>
							<div class='carousel-caption capa-alerta-1' style='background: !important;'>
								
								<span class='capa-inf-1'></span>
							</div>
						</a></div><div class='item '><a href='http://www.uca.edu.sv/seminariodemigracion/'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/03/banner-web-seminario-migraciones.jpg' alt=''  /></a> 
						<a href='http://www.uca.edu.sv/seminariodemigracion/'>
							<div class='carousel-caption capa-alerta-1' style='background: !important;'>
								
								<span class='capa-inf-1'></span>
							</div>
						</a></div><div class='item '><a href='http://www.uca.edu.sv/vida-estudiantil/'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/02/8.jpg' alt='Preinscripción e inscripción del Ciclo 01/2018'  /></a> 
						<a href='http://www.uca.edu.sv/vida-estudiantil/'>
							<div class='carousel-caption capa-alerta-1' style='background:#eb5218 !important;'>
								Preinscripción e inscripción del Ciclo 01/2018
								<span class='capa-inf-1'></span>
							</div>
						</a></div><div class='item '><a href='http://www.uca.edu.sv/acerca-de-la-uca/investigacion/'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/02/BANER-WEB-CONVOCATORIA-2018-FINANCIAMIENT-PROYECTS-INVESTIG-seleccionada.jpg' alt=''  /></a> 
						<a href='http://www.uca.edu.sv/acerca-de-la-uca/investigacion/'>
							<div class='carousel-caption capa-alerta-1' style='background: !important;'>
								
								<span class='capa-inf-1'></span>
							</div>
						</a></div></div><a class="left ant carousel-control" href="#banner" role="button" data-slide="prev" id="ant">
				<span class="glyphicon glyphicon-chevron-left" aria-hidden="true"></span>
				<span class="sr-only">Previous</span>
			</a>
			<a class="right sig carousel-control" href="#banner" role="button" data-slide="next" id="sig">
				<span class="glyphicon glyphicon-chevron-right" aria-hidden="true"></span>
				<span class="sr-only">Next</span>
			</a></div></div><div class="clearfix"></div><div class="separador-lg"></div></div></section><section>
<a name="eventos-noticias"></a>
	<div class="container xancla">
		<div class="col-md-12 text-center">
			<span class="titulo-apartado">
				<span class="fondo">
					Eventos<span class="hidden-xs"> y noticias
				</span>
			</span>
		</div>
		<div class="separador"></div>
		<div class="col-sm-6 col-md-5 cartelera-separador cartelera-portada">
			<div class="btn_x_right">
				<a href="http://www.uca.edu.sv/cartelera/" class="btn btn-primary">
					<span class="hidden-xs">Cartelera</span><span class="hidden-sm hidden-md hidden-lg">Más</span>
				</a>
			</div>
			<div class="separador"></div>
			
            <div class='cartelera'>
            <div class="fecha">
                <div class="dia">
                    18
                </div>
                <div class="mes">
                    MAR
                </div>
            </div>
        
            <div class="informacion">
                        <div class="clearfix"></div>
                        <div class="item_sub">                        
                            <a href="http://www.uca.edu.sv/cartelera/concierto-entre-rutilio-y-romero/">Concierto: Entre Rutilio y Romero, <em>Misa popular salvadoreña</em></a>                        
                            <div class="clearfix"></div>
                             
                            <div class="clearfix"></div>                        
                            <div class="separador"></div>
                        </div> 
                    
            </div>
            <div class="clearfix"></div>
        </div>
            <div class="clearfix"></div>
            <div class="separador"></div>
            <div class='cartelera cartelera-no-border'>
            <div class="fecha">
                <div class="dia">
                    21
                </div>
                <div class="mes">
                    MAR
                </div>
            </div>
        
            <div class="informacion">
                        <div class="clearfix"></div>
                        <div class="item_sub">                        
                            <a href="http://www.uca.edu.sv/cartelera/catedra-inaugural-licenciatura-en-comunicacion-social/">Cátedra inaugural del Ciclo 01/2018 de la Licenciatura en Comunicación Social</a>                        
                            <div class="clearfix"></div>
                             
                            <div class="clearfix"></div>                        
                            <div class="separador"></div>
                        </div> 
                    
            </div>
            <div class="clearfix"></div>
        </div>
            <div class="clearfix"></div>
            <div class="separador"></div>
            <div class='cartelera'>
            <div class="fecha">
                <div class="dia">
                    22
                </div>
                <div class="mes">
                    MAR
                </div>
            </div>
        
            <div class="informacion">
                        <div class="clearfix"></div>
                        <div class="item_sub">                        
                            <a href="http://www.uca.edu.sv/cartelera/presentacion-estudio-institucionalidad-del-agua/">Presentación del estudio <em>Institucionalidad del agua en América Latina</em></a>                        
                            <div class="clearfix"></div>
                             
                            <div class="clearfix"></div>                        
                            <div class="separador"></div>
                        </div> 
                    
            </div>
            <div class="clearfix"></div>
        </div>
            <div class="clearfix"></div>
            <div class="separador"></div>
			
		</div>
		<div class="separador hidden-sm hidden-md hidden-lg"></div>
		<div class="col-sm-6 col-md-4 hidden-sm hidden-md hidden-lg text-center">

			<span class="titulo-apartado">
				<span class="fondo">
					Noticias
				</span>
			</span>
		</div>
		<div class="separador hidden-sm hidden-md hidden-lg"></div>
		<div class="col-sm-6 col-md-4">
		<div class="btn_x_right">
				<a href="http://www.uca.edu.sv/noticias/" target="n_ventana" class="btn btn-primary">
					<span class="hidden-xs">Noticias UCA</span><span class="hidden-sm hidden-md hidden-lg">Más</span>
				</a>
			</div>
			<div class="separador"></div>
			                                
            <img src='/upload_w/8/archivo/1520892813-5aa6fb8dd2db5.jpg'  class='img-responsive'/>
            
                           
            <a href="http://uca.edu.sv/noticias/texto-5319">
                Por Carla Ayala
            </a><br />             
            <span class="color-2 fuente-14">12/03/2018</span>           
            <div class="clearfix"></div>
            <div class="separador hidden-sm hidden-md hidden-lg"></div>
        
		</div>
		<div class="col-sm-6 col-md-3 noticia-portada">
			

			<div class="separador hidden-xs"></div>
			<div class="separador hidden-xs"></div>

			                                
            
            <span class='fuente-16'>Editorial</span><br />
                           
            <a href="http://uca.edu.sv/noticias/texto-5331">
                &iquest;Otro mundo es posible?
            </a><br />             
            <span class="color-2 fuente-14">16/03/2018</span>           
            <div class="clearfix"></div>
            <div class="separador hidden-sm hidden-md hidden-lg"></div>
        

			<div class="separador hidden-xs"></div>
			<div class="separador hidden-xs"></div>
			                                
            
            <span class='fuente-16'>Opini&oacute;n</span><br />
                           
            <a href="http://uca.edu.sv/noticias/texto-5330">
                Desplante ciudadano
            </a><br />             
            <span class="color-2 fuente-14">15/03/2018</span>           
            <div class="clearfix"></div>
            <div class="separador hidden-sm hidden-md hidden-lg"></div>
        			
			
			
		</div>
	</div>
	
	<div class="separador hidden-sm hidden-md hidden-lg"></div>
</section><section>
<a name="lo-mas-reciente"></a>
		<div class="separador-lg hidden-xs "></div>
	<div class="container xancla">
		<div class="col-md-12 text-center">
		
			<span class="titulo-apartado">
				<span class="fondo">
					Lo más reciente
				</span>
			</span>
		</div>
		<div class="col-md-12 tabs-portada">		
			
		    <div class="separador"></div>			
			<ul class="nav nav-tabs nav-align responsive-tabs hidden-xs hidden-sm" role="tablist">
				<li role="presentation" class="active"><a href="#msj1" aria-controls="1" role="tab" data-toggle="tab" >Prácticas jurídicas</a></li><li role="presentation" ><a href="#msj2" aria-controls="2" role="tab" data-toggle="tab" >Informe de derechos humanos</a></li><li role="presentation" ><a href="#msj3" aria-controls="3" role="tab" data-toggle="tab" >Estudio socioeconómico 2017</a></li>				
			</ul>			
			<div class="tab-content cj-tab-content hidden-xs hidden-sm">
				<div class="separador"></div>
				<div role="tabpanel" class="tab-pane  in active" id="msj1"><p><img class="alignleft size-full wp-image-4241" src="http://www.uca.edu.sv/wp-content/uploads/2018/01/practicas-juridicas-lo-mas-reciente.jpg" alt="" width="500" height="182" />Dirigido a estudiantes, egresados y graduados de la Licenciatura en Ciencias Jurídicas de la UCA.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-dEhxus">Más información</a></p>
<p>&nbsp;</p></div><div role="tabpanel" class="tab-pane  " id="msj2"><p><img class="alignleft size-full wp-image-4107" src="http://www.uca.edu.sv/wp-content/uploads/2018/02/notificacion-informe-derechos-humanos.jpg" alt="" width="500" height="182" />El Instituto de Derechos Humanos de la UCA (Idhuca) presentó el informe “Balance de derechos humanos 2017”, que da cuenta de las violaciones a los derechos básicos, económicos y sociales, y valora el trabajo del sistema judicial.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-JZSCpY">Informe</a></p></div><div role="tabpanel" class="tab-pane  " id="msj3"><p><img class="size-full wp-image-4102 alignleft" src="http://www.uca.edu.sv/wp-content/uploads/2018/02/notificacion-analisis-socioeconomico.jpg" alt="" width="492" height="174" />Resultados del estudio “Análisis socioeconómico de El Salvador, año 2017”, elaborado por el Departamento de Economía. Entre los temas analizados destacan el mercado laboral y la fuerza de trabajo; la evolución de la productividad en El Salvador; demografía y desarrollo; desigualdad y polarización; política de ingreso; y política fiscal.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-hdSBuG">Estudio</a></p></div>			
			</div>		
		    
            <div class="panel-group hidden-md hidden-lg" id="accordion">
                
                    <div class="panel panel-default">
                        <a role="button" data-toggle="collapse" data-parent="#accordion" href="#collapse1">
                        <div class="panel-heading" >
                            <h4 class="panel-title">                                
                                Prácticas jurídicas                               
                            </h4>
                        </div>
                        </a>
                        <div id="collapse1" class="panel-collapse collapse   in">
                            <div class="panel-body">
                                <p><img class="alignleft size-full wp-image-4241" src="http://www.uca.edu.sv/wp-content/uploads/2018/01/practicas-juridicas-lo-mas-reciente.jpg" alt="" width="500" height="182" />Dirigido a estudiantes, egresados y graduados de la Licenciatura en Ciencias Jurídicas de la UCA.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-dEhxus">Más información</a></p>
<p>&nbsp;</p>
                            </div>
                        </div>
                    </div>
                    <div class="panel panel-default">
                        <a role="button" data-toggle="collapse" data-parent="#accordion" href="#collapse2">
                        <div class="panel-heading" >
                            <h4 class="panel-title">                                
                                Informe de derechos humanos                               
                            </h4>
                        </div>
                        </a>
                        <div id="collapse2" class="panel-collapse collapse ">
                            <div class="panel-body">
                                <p><img class="alignleft size-full wp-image-4107" src="http://www.uca.edu.sv/wp-content/uploads/2018/02/notificacion-informe-derechos-humanos.jpg" alt="" width="500" height="182" />El Instituto de Derechos Humanos de la UCA (Idhuca) presentó el informe “Balance de derechos humanos 2017”, que da cuenta de las violaciones a los derechos básicos, económicos y sociales, y valora el trabajo del sistema judicial.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-JZSCpY">Informe</a></p>
                            </div>
                        </div>
                    </div>
                    <div class="panel panel-default">
                        <a role="button" data-toggle="collapse" data-parent="#accordion" href="#collapse3">
                        <div class="panel-heading" >
                            <h4 class="panel-title">                                
                                Estudio socioeconómico 2017                               
                            </h4>
                        </div>
                        </a>
                        <div id="collapse3" class="panel-collapse collapse ">
                            <div class="panel-body">
                                <p><img class="size-full wp-image-4102 alignleft" src="http://www.uca.edu.sv/wp-content/uploads/2018/02/notificacion-analisis-socioeconomico.jpg" alt="" width="492" height="174" />Resultados del estudio “Análisis socioeconómico de El Salvador, año 2017”, elaborado por el Departamento de Economía. Entre los temas analizados destacan el mercado laboral y la fuerza de trabajo; la evolución de la productividad en El Salvador; demografía y desarrollo; desigualdad y polarización; política de ingreso; y política fiscal.</p>
<p style="text-align: center;"><a class="btn btn-primary" href="http://www.uca.edu.sv/-hdSBuG">Estudio</a></p>
                            </div>
                        </div>
                    </div>
            </div>
		</div>
	</div>
	<div class="separador-lg"></div>
</section><section>
<a name="orgullo-uca"></a>
	<div class="container xancla">
		<div class="separador-lg hidden-xs"></div>
		<div class="col-md-12 text-center">
		
			<span class="titulo-apartado">
				<span class="fondo">
					#OrgulloUCA
				</span>
			</span>
		</div>
		<div class="separador"></div>
	</div>
	<div class="container-fluid">		
		
		<div class="container-fluid hidden-sm hidden-md hidden-lg">
			<div class="col-md-12 no-padding">
			<div class="panel-group " id="accordion" role="tablist" aria-multiselectable="true">
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca1" aria-expanded="false" aria-controls="org_uca1">
					<div class="panel-heading" role="tab" id="heading_uca1">
						<h4 class="panel-title">
							
								David Barba aprobó con nota máxima su tesis de maestría en la UNAM
							
						</h4>
					</div>
					</a>

					<div id="org_uca1" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca1">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2018/02/David-Barba-web-700x535.jpg" class="img-responsive" />
							<p>David Barba, graduado de Ingeniería Civil, aprobó con nota máxima, 10, su tesis de la Maestría en Ingeniería Civil, con especialidad en Geotécnica, en la Universidad Nacional Autónoma de México. “Mi tema de tesis fue ‘Estudio del comportamiento de estructuras termoactivas, con énfasis en pilotes de energía’. Mi trabajo se enfocó en analizar su comportamiento desde el punto de vista geotécnico, evaluando los efectos que los cambios de temperatura tienen en el comportamiento mecánico de la cimentación. Pienso en posibles aportes de esta tecnología en El Salvador”.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca2" aria-expanded="false" aria-controls="org_uca2">
					<div class="panel-heading" role="tab" id="heading_uca2">
						<h4 class="panel-title">
							
								Ing. Erick Ramos en X Congreso Mundial de Ingeniería Química (España)
							
						</h4>
					</div>
					</a>

					<div id="org_uca2" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca2">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2018/02/Erick-Ramos-700x524.jpg" class="img-responsive" />
							<p>El ingeniero Erick Ramos, catedrático e investigador del Departamento de Ingeniería de Procesos y Ciencias Ambientales, participó en octubre de 2017 en el X Congreso Mundial de Ingeniería Química (Barcelona, España). Ramos, el único salvadoreño en el Congreso, expuso su investigación sobre el ácido anacárdico, un antioxidante natural, extraído de la cáscara de la nuez del marañón, que puede tener múltiples aplicaciones industriales y farmacéuticas, pero cuyo costo actual de producción es elevado. “Mi investigación plantea una forma más económica de extraer el ácido anacárdico".</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca3" aria-expanded="false" aria-controls="org_uca3">
					<div class="panel-heading" role="tab" id="heading_uca3">
						<h4 class="panel-title">
							
								Catalina Vásquez recibe reconocimiento en Chile
							
						</h4>
					</div>
					</a>

					<div id="org_uca3" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca3">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/12/Catalina-Vásquez-web-700x513.jpg" class="img-responsive" />
							<p>El 29 de noviembre de 2017, Catalina Vásquez, graduada de la Licenciatura en Comunicación Social, recibió de manos de la presidenta chilena, Michelle Bachelet, un reconocimiento por haber obtenido el mejor promedio (6.4 de 7.0) de entre los salvadoreños becados que estudian un posgrado en el país suramericano. “Crecimiento académico, profesional, pero sobre todo crecimiento personal”, así define Catalina su experiencia estudiando la Maestría en Ciencia Política en Chile, gracias a una beca a la que se hizo acreedora en 2016.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca4" aria-expanded="false" aria-controls="org_uca4">
					<div class="panel-heading" role="tab" id="heading_uca4">
						<h4 class="panel-title">
							
								Catedráticos DOE ganan primer lugar en concurso Conacyt 2017
							
						</h4>
					</div>
					</a>

					<div id="org_uca4" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca4">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/11/Ecomateriales-web-700x513.jpg" class="img-responsive" />
							<p>La investigación “Eco-materiales”, dirigida por los arquitectos Lizeth Rodríguez y Arturo Cisneros, catedráticos del Departamento de Organización del Espacio, ganó el primer lugar de la categoría Medio Ambiente del Premio Nacional en Investigación Científica y/o Tecnológica para Educación Superior y Centros de Investigación 2017, otorgado por el Viceministerio de Ciencia y Tecnología a través del Conacyt. “Ha sido un esfuerzo multi e interdisciplinario en el que han hecho sinergia académicos y estudiantes de la UCA”.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca5" aria-expanded="false" aria-controls="org_uca5">
					<div class="panel-heading" role="tab" id="heading_uca5">
						<h4 class="panel-title">
							
								Josué Arana, primer lugar en concurso iberoamericano
							
						</h4>
					</div>
					</a>

					<div id="org_uca5" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca5">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/11/josue-arana-700x506.jpg" class="img-responsive" />
							<p><span id="fbPhotoSnowliftCaption" class="fbPhotosPhotoCaption" tabindex="0" data-ft="{&quot;tn&quot;:&quot;K&quot;}"><span class="hasCaption">Josué Arana, egresado de Arquitectura de la UCA, ganó el primer lugar del Premio Vivir en Concreto, en el que participaron estudiantes de 35 universidades de 12 países de Iberoamérica y el Caribe. <br /> "La buena arquitectura, siempre nos lo han dicho acá [en la UCA],<span class="text_exposed_show"> va más allá. Me emocioné al crear esta vivienda, porque la pienso como si yo fuera a vivir ahí. No porque es para gente de escasos recursos voy a limitar el diseño; la idea es que puedan tener algo que valga la pena”.<br /> </span></span></span></p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca6" aria-expanded="false" aria-controls="org_uca6">
					<div class="panel-heading" role="tab" id="heading_uca6">
						<h4 class="panel-title">
							
								Obturador Libre gana primer lugar en Premio Pixels 2017
							
						</h4>
					</div>
					</a>

					<div id="org_uca6" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca6">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/12/obturadorlibre-700x517.jpg" class="img-responsive" />
							<p>Roberto Villalta, estudiante de Ingeniería Eléctrica, y Silsa Pineda, Laura Mejía y Luis Alvarado, de Comunicación Social, ganaron el primer lugar por Mejor Guion Original y Mejor Corto de Drama con su producción <em>El amor en tiempos del ciclo</em>, con la cual participaron en la categoría Tradicional del Premio Pixels 2017, entregado por la Dirección de Innovación y Calidad del Ministerio de Economía. Los jóvenes crearon la productora Obturador Libre, que les permite poner en práctica sus conocimientos académicos y ganar experiencia en el ámbito profesional.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca7" aria-expanded="false" aria-controls="org_uca7">
					<div class="panel-heading" role="tab" id="heading_uca7">
						<h4 class="panel-title">
							
								María Eugenia Gálvez en Lituania
							
						</h4>
					</div>
					</a>

					<div id="org_uca7" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca7">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/09/21551855_10155862952932722_414412634320802076_o-700x394.jpg" class="img-responsive" />
							<p>María Eugenia Gálvez, de la Licenciatura en Mercadeo, cursó un semestre en la Universidad de Vilnius (Lituania), tras obtener una beca otorgada por el Programa Erasmus Plus, de la Unión Europea. “Hay que quitarse el miedo de fracasar y dejar de minimizar las cosas que hacemos. En El Salvador, todo está polarizado, no hay disposición de ponerse en el lugar del otro. Afuera uno entiende lo necesario que es tener empatía para progresar”, afirma.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca8" aria-expanded="false" aria-controls="org_uca8">
					<div class="panel-heading" role="tab" id="heading_uca8">
						<h4 class="panel-title">
							
								P. José María Tojeira recibe premio CLACSO 50 años
							
						</h4>
					</div>
					</a>

					<div id="org_uca8" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca8">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/11/jose-maria-tojeira-orgullouca-700x506.jpg" class="img-responsive" />
							<p>Por sus aportes a la defensa y promoción de los derechos humanos, su compromiso con las víctimas de la violencia y su lucha a favor de los sectores populares, el padre José María Tojeira, director del Idhuca, recibió el premio CLACSO 50 años. “Acepto su distinción como un homenaje comprometedor con todos aquellos que a lo largo de estos años difíciles nos han mostrado el camino de la generosidad social y la inteligencia creativa”, dijo el P. Tojeira en su mensaje a CLACSO.</p>
						</div>
					</div>
				</div>


				
				
			


				<div class="panel panel-default">
				<a class="collapsed" role="button" data-toggle="collapse" data-parent="#accordion" href="#org_uca9" aria-expanded="false" aria-controls="org_uca9">
					<div class="panel-heading" role="tab" id="heading_uca9">
						<h4 class="panel-title">
							
								Nelson Quintanilla rumbo a Canadá
							
						</h4>
					</div>
					</a>

					<div id="org_uca9" class="panel-collapse collapse" role="tabpanel" aria-labelledby="heading_uca9">
						<div class="panel-body">
							<img  src="http://www.uca.edu.sv/wp-content/uploads/2017/09/21317411_10155821226647722_2056020686704873104_n-700x531.jpg" class="img-responsive" />
							<p>Nelson Quintanilla tiene 22 años, cursa cuarto año de Ingeniería Eléctrica y es beneficiario del Programa de Becas Parciales UCA. . Gracias a su buen desempeño académico, obtuvo una beca de intercambio, otorgada por el Programa Líderes Emergentes de las Américas, que le permitirá estudiar un semestre en la Universidad de New Brunswick (Canadá). Durante su estadía en Canadá, cursará materias como Ingeniería Económica, Introducción a la Mecatrónica, Leyes y Ética para Ingeniería, y Cambio Climático y Ciudad.</p>
						</div>
					</div>
				</div>


				
				
			</div>
			</div>
		</div>



	<div class="container-fluid no-padding hidden-xs">
		<div class="col-md-12 no-padding">
			<div id="orgulloUCA" class="carousel slide" data-ride="carousel"><div class="carousel-inner anim" role="listbox"><div class='item active'><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/02/David-Barba-web-700x535.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>David Barba, graduado de Ingeniería Civil, aprobó con nota máxima, 10, su tesis de la Maestría en Ingeniería Civil, con especialidad en Geotécnica, en la Universidad Nacional Autónoma de México. “Mi tema de tesis fue ‘Estudio del comportamiento de estructuras termoactivas, con énfasis en pilotes de energía’. Mi trabajo se enfocó en analizar su comportamiento desde el punto de vista geotécnico, evaluando los efectos que los cambios de temperatura tienen en el comportamiento mecánico de la cimentación. Pienso en posibles aportes de esta tecnología en El Salvador”.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2018/02/Erick-Ramos-700x524.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>El ingeniero Erick Ramos, catedrático e investigador del Departamento de Ingeniería de Procesos y Ciencias Ambientales, participó en octubre de 2017 en el X Congreso Mundial de Ingeniería Química (Barcelona, España). Ramos, el único salvadoreño en el Congreso, expuso su investigación sobre el ácido anacárdico, un antioxidante natural, extraído de la cáscara de la nuez del marañón, que puede tener múltiples aplicaciones industriales y farmacéuticas, pero cuyo costo actual de producción es elevado. “Mi investigación plantea una forma más económica de extraer el ácido anacárdico".</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/12/Catalina-Vásquez-web-700x513.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>El 29 de noviembre de 2017, Catalina Vásquez, graduada de la Licenciatura en Comunicación Social, recibió de manos de la presidenta chilena, Michelle Bachelet, un reconocimiento por haber obtenido el mejor promedio (6.4 de 7.0) de entre los salvadoreños becados que estudian un posgrado en el país suramericano. “Crecimiento académico, profesional, pero sobre todo crecimiento personal”, así define Catalina su experiencia estudiando la Maestría en Ciencia Política en Chile, gracias a una beca a la que se hizo acreedora en 2016.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/11/Ecomateriales-web-700x513.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>La investigación “Eco-materiales”, dirigida por los arquitectos Lizeth Rodríguez y Arturo Cisneros, catedráticos del Departamento de Organización del Espacio, ganó el primer lugar de la categoría Medio Ambiente del Premio Nacional en Investigación Científica y/o Tecnológica para Educación Superior y Centros de Investigación 2017, otorgado por el Viceministerio de Ciencia y Tecnología a través del Conacyt. “Ha sido un esfuerzo multi e interdisciplinario en el que han hecho sinergia académicos y estudiantes de la UCA”.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/11/josue-arana-700x506.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p><span id="fbPhotoSnowliftCaption" class="fbPhotosPhotoCaption" tabindex="0" data-ft="{&quot;tn&quot;:&quot;K&quot;}"><span class="hasCaption">Josué Arana, egresado de Arquitectura de la UCA, ganó el primer lugar del Premio Vivir en Concreto, en el que participaron estudiantes de 35 universidades de 12 países de Iberoamérica y el Caribe. <br /> "La buena arquitectura, siempre nos lo han dicho acá [en la UCA],<span class="text_exposed_show"> va más allá. Me emocioné al crear esta vivienda, porque la pienso como si yo fuera a vivir ahí. No porque es para gente de escasos recursos voy a limitar el diseño; la idea es que puedan tener algo que valga la pena”.<br /> </span></span></span></p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/12/obturadorlibre-700x517.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>Roberto Villalta, estudiante de Ingeniería Eléctrica, y Silsa Pineda, Laura Mejía y Luis Alvarado, de Comunicación Social, ganaron el primer lugar por Mejor Guion Original y Mejor Corto de Drama con su producción <em>El amor en tiempos del ciclo</em>, con la cual participaron en la categoría Tradicional del Premio Pixels 2017, entregado por la Dirección de Innovación y Calidad del Ministerio de Economía. Los jóvenes crearon la productora Obturador Libre, que les permite poner en práctica sus conocimientos académicos y ganar experiencia en el ámbito profesional.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/09/21551855_10155862952932722_414412634320802076_o-700x394.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>María Eugenia Gálvez, de la Licenciatura en Mercadeo, cursó un semestre en la Universidad de Vilnius (Lituania), tras obtener una beca otorgada por el Programa Erasmus Plus, de la Unión Europea. “Hay que quitarse el miedo de fracasar y dejar de minimizar las cosas que hacemos. En El Salvador, todo está polarizado, no hay disposición de ponerse en el lugar del otro. Afuera uno entiende lo necesario que es tener empatía para progresar”, afirma.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/11/jose-maria-tojeira-orgullouca-700x506.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>Por sus aportes a la defensa y promoción de los derechos humanos, su compromiso con las víctimas de la violencia y su lucha a favor de los sectores populares, el padre José María Tojeira, director del Idhuca, recibió el premio CLACSO 50 años. “Acepto su distinción como un homenaje comprometedor con todos aquellos que a lo largo de estos años difíciles nos han mostrado el camino de la generosidad social y la inteligencia creativa”, dijo el P. Tojeira en su mensaje a CLACSO.</p></div></div></div></div><div class='item '><div class='container'><div class='col-md-5'><img  src='http://www.uca.edu.sv/wp-content/uploads/2017/09/21317411_10155821226647722_2056020686704873104_n-700x531.jpg'' class='img-responsive' /></div><div class='col-md-7 text-center'>
				<div class='vcenter div335min fuente-24'><p>Nelson Quintanilla tiene 22 años, cursa cuarto año de Ingeniería Eléctrica y es beneficiario del Programa de Becas Parciales UCA. . Gracias a su buen desempeño académico, obtuvo una beca de intercambio, otorgada por el Programa Líderes Emergentes de las Américas, que le permitirá estudiar un semestre en la Universidad de New Brunswick (Canadá). Durante su estadía en Canadá, cursará materias como Ingeniería Económica, Introducción a la Mecatrónica, Leyes y Ética para Ingeniería, y Cambio Climático y Ciudad.</p></div></div></div></div></div><a class="left antt carousel-control" href="#orgulloUCA" role="button" data-slide="prev" id="ant">
			<span class="glyphicon glyphicon-chevron-left" aria-hidden="true"></span>
			<span class="sr-only">Previous</span>
		</a>
		<a class="right sigg carousel-control" href="#orgulloUCA" role="button" data-slide="next" id="sig">
			<span class="glyphicon glyphicon-chevron-right" aria-hidden="true"></span>
			<span class="sr-only">Next</span>
		</a></div></div><div class="clearfix"></div><div class="separador"></div></div>
	</div>
	<div class="separador-lg"></div>
</section><footer>
    <div class="separador"></div>
    <div class="separador"></div>
    <div class="container-fluid fondo-1">
        <div class="container">
            <div class="col-md-6 footer">
                <a href="http://www.facebook.com/UCA.ElSalvador"><img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/facebook.png" data-toggle="tooltip" data-placement="bottom" title="Síguenos en Facebook" /></a>
                <a href="http://twitter.com/UCA_ES"><img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/twitter.png" data-toggle="tooltip" data-placement="bottom" title="Síguenos en Twitter"/></a>
                <a href="https://www.instagram.com/uca_elsalvador/"><img src="http://www.uca.edu.sv/wp-content/themes/kubo/images/instagram.png" data-toggle="tooltip" data-placement="bottom" title="Síguenos en Instagram" /></a>
                <div class="clearfix"></div>
                            </div>
            <div class="col-md-6 footer text-right">
                <h3 class="no-margin">
                    Universidad Centroamericana José Simeón Cañas
                </h3>
                Bulevar Los Próceres, Antiguo Cuscatlán, La Libertad, El Salvador, Centroamérica <br />
                (503) 2210-6600 <a href="mailto:direccion.comunicaciones@uca.edu.sv">direccion.comunicaciones@uca.edu.sv</a>
                <div class="clearfix"></div>
            </div>
        </div>
    </div>
</footer>

<script src="https://ajax.googleapis.com/ajax/libs/jquery/1.12.4/jquery.min.js"></script>
<script src="http://www.uca.edu.sv/wp-content/themes/kubo/js/bootstrap.min.js"></script>

<script type="text/javascript">
    
$(document).ready(function(){
    var windowHeight = $(window).height();
    $(window).resize(function() {
        var windowHeight = $(window).height();
        $('.ancho').css('min-height',windowHeight-300);
    });

    urlHash = window.location.href;
    v_url= urlHash.indexOf( '#' );  

$('.menuG a').click(function(){
    $('.xancla').addClass('ancla_uca');
})
        var url = window.location.hash; //href;
        var hash = url.substring(url.indexOf("#")+1);
        
        if(url!==""){
            //$('.'+hash).addClass('ancla_uca');
            $('.xancla').addClass('ancla_uca');
               
                    //$('.'+hash).delay( 800 ).removeClass('ancla_uca');
            
            
        }

});
//$('.collapse').collapse();
</script>
<script src="http://www.uca.edu.sv/wp-content/themes/kubo/js/jquery.validate.min.js"></script>
<script src="http://www.uca.edu.sv/wp-content/themes/kubo/js/tema.js?697961078"></script>

<!-- Modal -->
<div class="modal fade" id="comunicaciones" tabindex="-1" role="dialog" aria-labelledby="contacto">
	<div class="modal-dialog" role="document">
		<div class="modal-content">
			<div class="modal-header">
				<button type="button" class="close" data-dismiss="modal" aria-label="Close"><span aria-hidden="true">&times;</span></button>
				<h4 class="modal-title" id="contacto">Buscar contenido</h4>
			</div>
			<div class="modal-body">
				<form action="http://www.uca.edu.sv/buscador/" method="get" id="form_bq">
                        <div class="input-group ">
                            <input type="text" class="form-control" placeholder="Buscar" name="q" id="q" value="">
                            <span class="input-group-btn" >
                                <button class="btn btn-default" type="submit"><span class="glyphicon glyphicon-search"></span></button>
                            </span>
                        </div>
                    </form>
			</div>
			<div class="modal-footer">
				<button type="button" class="btn btn-default" data-dismiss="modal">Cerrar</button>				
			</div>
		</div>
	</div>
</div>
</body>
</html>