<!DOCTYPE html>
<html lang="es-ES" prefix="og: http://ogp.me/ns#">
  
<head>
  <script async src="https://www.googletagmanager.com/gtag/js?id=UA-107318580-2"></script>
<script>
  window.dataLayer = window.dataLayer || [];
  function gtag(){dataLayer.push(arguments)};
  gtag('js', new Date());

  gtag('config', 'UA-107318580-2');
</script>
  
    <meta http-equiv="Content-Type" content="text/html; charset=UTF-8"/>

    <meta http-equiv="X-UA-Compatible" content="IE=Edge">

    <meta name="viewport" content="width=device-width, initial-scale=1, maximum-scale=1">

    <!-- For use in JS files -->
    <script type="text/javascript">
        var template_dir = "http://www.uees.edu.sv/wp-content/themes/invent5";
    </script>

    <link rel="profile" href="http://gmpg.org/xfn/11"/>

    <link rel="pingback" href="http://www.uees.edu.sv/xmlrpc.php"/>

    <script type="text/javascript">var mo_options = mo_options || {};mo_options.disable_back_to_top = false;mo_options.sticky_menu = true;mo_options.theme_skin = "#203864";mo_options.theme_directory_url = "http://www.uees.edu.sv/wp-content/themes/invent5";mo_options.slider_chosen="Revolution";mo_options.disable_smooth_page_load=false;mo_options.disable_animations_on_page=false;mo_options.disable_smooth_scroll=true;</script>
    <title>Inicio - Universidad Evangélica de El Salvador</title>

	<!-- Meta Tag Manager -->
	<meta name="description" content="Universidad Evangelica de El Salvador con Educación de Calidad y Valores Cristianos" />
	<meta name="keywords" content="Universidad, carreras, facultades, ingenierías, medicina, enfermería,administración de empresas, ciencias Jurídicas, ciencias Sociales,Computacion, redes, Ngocios, Mercadeo, Técnico, Recursos Humanos, Psicología,   Doctorado en Cirugía Dental, marketing, posgrados, pre grado, matricula, becas, nuevo ingreso, admisión , aranceles, Portal de Estudiante, portal del docente, proyección social, graduados , biblioteca UEES, uees,cooperación Internacional, publicaciones, deportes,arte y cultura, memoria de labores, beneficios, orientación vocacional, secretaria de Asuntos Espirituales, admisión de extranjeros, preguntas frecuentes, calendario académico, campus virtual uees" />
	<!-- / Meta Tag Manager -->

<!-- This site is optimized with the Yoast SEO plugin v6.2 - https://yoa.st/1yg?utm_content=6.2 -->
<link rel="canonical" href="http://www.uees.edu.sv/" />
<meta property="og:locale" content="es_ES" />
<meta property="og:type" content="website" />
<meta property="og:title" content="Inicio - Universidad Evangélica de El Salvador" />
<meta property="og:description" content="Bienvenidos a la Universidad Evangélica de El Salvador MensajesCatálogo InstitucionalModelo EducativoConveniosMensaje de BienvenidaEstimados Estudiantes:Las bases filosóficas y pedagógicas de nuestro proyecto educativo nos han orientado desde la fundación de la Universidad en 1981, a asumir los retos y compromisos de la Educación Superior en El Salvador. Esto significa para nosotros el reconocimiento de la importancia &hellip;" />
<meta property="og:url" content="http://www.uees.edu.sv/" />
<meta property="og:site_name" content="Universidad Evangélica de El Salvador" />
<meta property="og:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio3.png" />
<meta property="og:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio44-1.png" />
<meta property="og:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio1.png" />
<meta property="og:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio2.png" />
<meta property="og:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logopanalExok.png" />
<meta name="twitter:card" content="summary_large_image" />
<meta name="twitter:description" content="Bienvenidos a la Universidad Evangélica de El Salvador MensajesCatálogo InstitucionalModelo EducativoConveniosMensaje de BienvenidaEstimados Estudiantes:Las bases filosóficas y pedagógicas de nuestro proyecto educativo nos han orientado desde la fundación de la Universidad en 1981, a asumir los retos y compromisos de la Educación Superior en El Salvador. Esto significa para nosotros el reconocimiento de la importancia [&hellip;]" />
<meta name="twitter:title" content="Inicio - Universidad Evangélica de El Salvador" />
<meta name="twitter:site" content="@ueesoficial" />
<meta name="twitter:image" content="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio3.png" />
<meta name="twitter:creator" content="@ueesoficial" />
<script type='application/ld+json'>{"@context":"http:\/\/schema.org","@type":"WebSite","@id":"#website","url":"http:\/\/www.uees.edu.sv\/","name":"Universidad Evang\u00e9lica de EL Salvador","alternateName":"UEES, universidad evangelica de El Salvador, Escuela de posgrado, facultades, carreras, estudios,","potentialAction":{"@type":"SearchAction","target":"http:\/\/www.uees.edu.sv\/?s={search_term_string}","query-input":"required name=search_term_string"}}</script>
<script type='application/ld+json'>{"@context":"http:\/\/schema.org","@type":"Organization","url":"http:\/\/www.uees.edu.sv\/","sameAs":["https:\/\/www.facebook.com\/ueesoficial\/","https:\/\/www.instagram.com\/explore\/locations\/1012393993\/","https:\/\/www.youtube.com\/channel\/UCZ3m1ZKVzbsyuB3ZZlgXegA","https:\/\/twitter.com\/ueesoficial"],"@id":"#organization","name":"Universidad Evang\u00e9lica de EL Salvador","logo":"http:\/\/www.uees.edu.sv\/wp-content\/uploads\/2017\/06\/logouees.png"}</script>
<meta name="google-site-verification" content="mV_xAokPQauX2PQZg_acuUfbyycvc6trZtIOiBak2BI" />
<!-- / Yoast SEO plugin. -->

<link rel='dns-prefetch' href='//html5shiv.googlecode.com' />
<link rel='dns-prefetch' href='//s.w.org' />
<link rel="alternate" type="application/rss+xml" title="Universidad Evangélica de El Salvador &raquo; Feed" href="http://www.uees.edu.sv/?feed=rss2" />
<link rel="alternate" type="application/rss+xml" title="Universidad Evangélica de El Salvador &raquo; RSS de los comentarios" href="http://www.uees.edu.sv/?feed=comments-rss2" />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/www.uees.edu.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.7.5"}};
			!function(a,b,c){function d(a){var b,c,d,e,f=String.fromCharCode;if(!k||!k.fillText)return!1;switch(k.clearRect(0,0,j.width,j.height),k.textBaseline="top",k.font="600 32px Arial",a){case"flag":return k.fillText(f(55356,56826,55356,56819),0,0),!(j.toDataURL().length<3e3)&&(k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,65039,8205,55356,57096),0,0),b=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,55356,57096),0,0),c=j.toDataURL(),b!==c);case"emoji4":return k.fillText(f(55357,56425,55356,57341,8205,55357,56507),0,0),d=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55357,56425,55356,57341,55357,56507),0,0),e=j.toDataURL(),d!==e}return!1}function e(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var f,g,h,i,j=b.createElement("canvas"),k=j.getContext&&j.getContext("2d");for(i=Array("flag","emoji4"),c.supports={everything:!0,everythingExceptFlag:!0},h=0;h<i.length;h++)c.supports[i[h]]=d(i[h]),c.supports.everything=c.supports.everything&&c.supports[i[h]],"flag"!==i[h]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[i[h]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(g=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",g,!1),a.addEventListener("load",g,!1)):(a.attachEvent("onload",g),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),f=c.source||{},f.concatemoji?e(f.concatemoji):f.wpemoji&&f.twemoji&&(e(f.twemoji),e(f.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='stylesheet' id='formidable-css'  href='http://www.uees.edu.sv/wp-content/plugins/formidable/css/formidableforms.css?ver=382242' type='text/css' media='all' />
<link rel='stylesheet' id='flowplayer-css-css'  href='http://www.uees.edu.sv/wp-content/plugins/easy-video-player/lib/skin/skin.css?ver=4.7.5' type='text/css' media='all' />
<link rel='stylesheet' id='lsow-frontend-styles-css'  href='http://www.uees.edu.sv/wp-content/plugins/livemesh-siteorigin-widgets/assets/css/lsow-frontend.css?ver=1.7.3' type='text/css' media='all' />
<link rel='stylesheet' id='lsow-icomoon-styles-css'  href='http://www.uees.edu.sv/wp-content/plugins/livemesh-siteorigin-widgets/assets/css/icomoon.css?ver=1.7.3' type='text/css' media='all' />
<link rel='stylesheet' id='tp_twitter_plugin_css-css'  href='http://www.uees.edu.sv/wp-content/plugins/recent-tweets-widget/tp_twitter_plugin.css?ver=1.0' type='text/css' media='screen' />
<link rel='stylesheet' id='rs-plugin-settings-css'  href='http://www.uees.edu.sv/wp-content/plugins/revslider/public/assets/css/settings.css?ver=5.4.1' type='text/css' media='all' />
<style id='rs-plugin-settings-inline-css' type='text/css'>
#rs-demo-id {}
</style>
<link rel='stylesheet' id='siteorigin-panels-front-css'  href='http://www.uees.edu.sv/wp-content/plugins/siteorigin-panels/css/front-flex.min.css?ver=2.6.3' type='text/css' media='all' />
<link rel='stylesheet' id='sow-image-default-642c5433d908-css'  href='http://www.uees.edu.sv/wp-content/uploads/siteorigin-widgets/sow-image-default-642c5433d908.css?ver=4.7.5' type='text/css' media='all' />
<link rel='stylesheet' id='megamenu-css'  href='http://www.uees.edu.sv/wp-content/uploads/maxmegamenu/style.css?ver=a8fdde' type='text/css' media='all' />
<link rel='stylesheet' id='dashicons-css'  href='http://www.uees.edu.sv/wp-includes/css/dashicons.min.css?ver=4.7.5' type='text/css' media='all' />
<link rel='stylesheet' id='pretty-photo-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/prettyPhoto.css?ver=4.7.5' type='text/css' media='screen' />
<link rel='stylesheet' id='icon-fonts-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/icon-fonts.css?ver=4.7.5' type='text/css' media='screen' />
<link rel='stylesheet' id='style-theme-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/style.css?ver=4.7.5' type='text/css' media='all' />
<!--[if IE 8]>
<link rel='stylesheet' id='style-ie8-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/ie8.css?ver=4.7.5' type='text/css' media='screen' />
<![endif]-->
<!--[if IE 9]>
<link rel='stylesheet' id='style-ie9-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/ie9.css?ver=4.7.5' type='text/css' media='screen' />
<![endif]-->
<link rel='stylesheet' id='animate-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/animate.css?ver=4.7.5' type='text/css' media='screen' />
<link rel='stylesheet' id='js_composer_front-css'  href='http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/css/js_composer.min.css?ver=5.2' type='text/css' media='all' />
<link rel='stylesheet' id='style-plugins-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/css/plugins.css?ver=4.7.5' type='text/css' media='all' />
<link rel='stylesheet' id='style-custom-css'  href='http://www.uees.edu.sv/wp-content/themes/invent5/custom/custom.css?ver=4.7.5' type='text/css' media='all' />
<style id='style-custom-inline-css' type='text/css'>
@import url("//fonts.googleapis.com/css?family=Lato");

h1,h2,h3,h4,h5,h6, .slogan1, #slider-area .flex-caption a, ul.tab-list li a, ul.member-list li a, .number-stats .number-stat .number, #mobile-menu .menu-header, .heading2 .subtitle span, .video-section .video-header .header-content .text, .ytp-video-section .video-header .header-content .text, .single .number-stats .number-stat .number, #content .marketing-banner ol.simple-list a, #content .marketing-banner ol.events-list a, .course-details .header, .staff-details .header, .department-details .header, .department-details .contact-person .name, .post-snippets .hentry .entry-title, .post-snippets .type-course .img-wrap .type-info .post-title, .post-snippets .type-news .img-wrap .type-info .post-title, .post-snippets .type-staff .img-wrap .type-info .post-title, .post-snippets .type-department .img-wrap .type-info .post-title, .single-event .heading-title, .single-location .heading-title, .css-events-list .events-table td a, table.em-calendar thead .month_name, .tribe-events-venue-widget .tribe-venue-widget-venue .tribe-venue-widget-venue-name a, .tribe-events-countdown-widget div.tribe-countdown-text, .tribe-events-countdown-widget .tribe-countdown-number, .heading2 .title, .number-stats .number-stat .stats-title, .image-info .post-title, ul.post-list .entry-title a, #learndash_next_prev_link, #learndash_back_to_lesson {font-family:"H1, "Lato", Arial, Helvetica, Verdana, sans-serif";}
#learndash_lessons, #learndash_quizzes, .expand_collapse, .notavailable_message, #learndash_lesson_topics_list div > strong, #learndash_lesson_topics_list div ul > li .sn, .learndash_profile_heading, #learndash_profile a, #learndash_profile div {font-family:"H1, "Lato", Arial, Helvetica, Verdana, sans-serif" !important;}
h1,h2,h3,h4,h5,h6, .slogan1, .heading2 .title {letter-spacing:3px;}
body, button, .button, input[type=button], input[type="submit"], input[type="reset"], .timeline-footer .event-date, .timeline-footer .event-category, .subtitle, .client-testimonials2 .header cite, .page-links a, .page-links a:visited, .pagination a, .pagination a:visited, .pagination span.current, .post-snippets .type-course .course-id, .course-details .course-information .label, .dropdown-menu-wrap ul li a, blockquote .author, blockquote em, blockquote i, blockquote cite, #top-header-area ul.contact-info li, #top-header-area ul.contact-info li a, .comment-reply-link, .comment-edit-link, .comment-reply-link:visited, .comment-edit-link:visited, #course_navigation .learndash_nevigation_lesson_topics_list .lesson a, .widget_course_return, #course_navigation .widget_course_return a, #course_navigation .learndash_topic_widget_list a > span, #course_navigation .learndash_nevigation_lesson_topics_list .lesson, .widget_ldcourseinfo #ld_course_info #course_progress_details > strong, .widget_course_return, #course_navigation .widget_course_return a, .wpProQuiz_forms table td label, .wpProQuiz_maxtrixSortText, .wpProQuiz_sortable, .wpProQuiz_sortStringItem {font-family:"Arial";}
#learndash_lessons a, #learndash_quizzes a, .expand_collapse a, .learndash_topic_dots a, .learndash_topic_dots a > span, #learndash_lesson_topics_list span a, #learndash_profile a, #learndash_profile a span, .wpProQuiz_questionListItem input[type="radio"], .wpProQuiz_questionListItem input[type="checkbox"], .wpProQuiz_questionListItem span {font-family:"Arial" !important;}
cite, em, i, #author-widget .author-name, blockquote, .pullquote, .rss-block, ul.post-list .published, ul.post-list .byline, ul.post-list .entry-meta, .entry-meta span, .entry-meta span a, .comment-author cite, .comment-byline, #services-icon-list .sub, .post-snippets .byline {font-family:"Lato";}
body{font-size:15px;}
#header .inner .wrap {height:60px !important;}
#primary-menu > ul.menu > li > a {font-size:17px !important;}
#primary-menu ul.menu > li.sfHover > a, #primary-menu > ul.menu > li > a:hover { color:#f9e500 !important; }
.dropdown-menu-wrap ul.sub-menu { background-color: #ffffff;}
.dropdown-menu-wrap ul.sub-menu li { border: none;}
.dropdown-menu-wrap ul.sub-menu > li a { color:#000000 !important;font-size:16px !important;}
.dropdown-menu-wrap ul.sub-menu li:hover, .dropdown-menu-wrap ul.sub-menu li.sfHover { background-color: #000000}
.dropdown-menu-wrap ul.sub-menu li:hover a, .dropdown-menu-wrap ul.sub-menu li.sfHover a { color:#6d6d6d !important;}
#main {background-color:#ffffff;background-image: none;background-attachment: fixed;background-size: cover;}
#pricing-action .pointing-arrow img { opacity: 0 }
/* ============== START - Skin Styles ============= */

th { background: #203864; }

/* ------- The links --------- */
a, a:active, a:visited { color: #203864; }
a:hover { color: #888; }
.dark-bg a { color: #203864 !important; }

blockquote .author, blockquote em, blockquote i, blockquote cite { color: #203864; }

.dropdown-menu-wrap ul.sub-menu li:hover, .dropdown-menu-wrap ul.sub-menu li.sfHover { background: #203864; }
#primary-menu > ul.menu > li:hover > ul.sub-menu { border-color: #203864; }
#primary-menu .hover-bg { border-color: #203864;}
#title-area { background: #203864; }
#custom-title-area { background: #203864; }

.post-list .entry-title a:hover, .post-list .entry-title a:visited { color: #203864; }
.sticky .entry-snippet { border-color: #203864;}
.entry-terms.multi-color .news_category, .entry-terms.multi-color .category { background-color: #203864; }
a.more-link:hover { color: #203864; }
a.comment-reply-link, a.comment-edit-link { background-color: #203864; }
a.comment-reply-link:visited, a.comment-edit-link:visited { background-color: #203864; }
button, .button, input[type=button], input[type="submit"], input[type="reset"] { background-color: #203864; border-color: #203864;}
.button.theme:hover { background: #203864 !important; }
.button.theme { border-color: #203864 !important; }


.segment .flex-control-nav li a:hover, .segment .flex-control-nav li a.flex-active { background-color: #203864; }

#flickr-widget .flickr_badge_image img:hover { border-color: #203864; }
ul#recentcomments li.recentcomments a { color: #203864; }
.tagcloud a:hover { background-color: #203864; }
input#mc_signup_submit { background-color: #203864 !important; }

.header-fancy span { background-color: #203864; }
h3.fancy-header { background-color: #203864;}

.skill-bar-content { background: #203864; }
.slogan1 .highlight, .slogan1 .highlight h2 { color: #203864; }
.heading2 .subtitle span { color: #203864; }
.heading1.separator .title:after, .heading2.separator .title:after { background: #203864; }
h4.subheading:after, h3.subheading:after { border-color: #203864; }

.segment.slogan blockquote .footer cite { color: #203864; }
.portfolio-label { color: #203864; }
.portfolio-index i:hover { color: #203864; }
#showcase-filter a:hover, #showcase-filter a.active, #showcase-links a:hover, #showcase-links a.active { background: #203864; border-color: #203864; }

.stats-bar-content { background: #203864; }
.number-stats .number-stat .number { color: #203864;}
.number-stats .number-stat .icon-wrap { background: #203864; }

.pricing-table .pricing-plan.highlight .top-header { background-color: #203864; }
.pricing-table .plan-details ul li i { color: #203864; }

.testimonials2-slider-container blockquote cite i { background-color: #203864; }
.client-testimonials2 .header cite { color: #203864;}
#services-icon-list div.icon { color: #203864;}
#services-icon-list .sub { color: #203864;}
.features-list-alternate i { color: #203864; }
ul.member-list { border-color: #203864; }
ul.member-list li a.visible, ul.member-list li a.flex-active { border-color: #203864; }
ul.member-list li a:hover { color: #203864; }
#showcase-filter a:hover { background: #203864; border-color: #203864; }

.timeline-item:before { background: #203864; }
.timeline-footer .event-category i { color: #203864; }

.course-details .header, .staff-details .header, .department-details .header { background: #203864; }
.post-snippets .type-course .course-id { background: #203864; }



#column-shortcode-section p { background: #203864; }

.top-of-page a:hover, .post-list .byline a, .post-list .byline a:active, .post-list .byline a:visited,
#content .hentry h2.entry-title a:hover, .entry-meta span i, .read-more a, .loop-nav a:hover,
.sidebar li > a:hover, .sidebar li:hover > a, #sidebars-footer .widget_text a.small, #sidebars-footer .widget_text a.small:visited,
#home-intro h2 span, .team-member:hover h3 a, .post-snippets .hentry .entry-title a:hover { color: #203864; }

.widget.widget_nav_menu ul li.current_page_item > a { background: #203864; }

.bx-wrapper .bx-pager.bx-default-pager a:hover, .bx-wrapper .bx-pager.bx-default-pager a.active,
.page-links a, .page-links a:visited, .pagination a, .pagination a:visited,
.profile-header img:hover { background: #203864; }

#styleswitcher-button i { color: #203864 !important; }

.profile-header .socials { background: rgba(32, 56 , 100, 0.7);}
input:focus, textarea:focus, #content .contact-form input:focus, #content .contact-form textarea:focus,
#footer .contact-form input:focus, #footer .contact-form textarea:focus { border-color: rgba(32, 56 , 100, 0.8); }
#home2-heading .heading2 h2, #home3-heading .heading2 h2, .team-member .team-member-hover { background: rgba(32, 56 , 100, 0.7); }

#footer .button:hover, #footer button:hover, #footer input[type="button"]:hover, #footer input[type="submit"]:hover, #footer input[type="reset"]:hover {
background-color: #203864 !important;
border-color: #203864 !important;
}

.tabs .current, .tabs .current:hover, .tabs li.current a { border-top-color: #203864; }
.toggle-label:hover, .active-toggle .toggle-label:hover { background-color: #203864; }

ul.tab-list, ul.member-list { border-bottom: 1px solid #203864; }
ul.tab-list li a.visible, ul.tab-list li a.flex-active, ul.member-list li a.visible, ul.member-list li a.flex-active { border-bottom: 3px solid #203864; }
ul.tab-list li a:hover, ul.member-list li a:hover { color: #203864; }

.sidebar .text-content a, #footer .text-content a { color: #203864; }

.gallery-carousel .carousel-container .owl-carousel.owl-theme .owl-prev, .gallery-carousel .carousel-container .owl-carousel.owl-theme .owl-next { background: #203864; }

/* Plugins Skins Styles */

/*---------- Events Manager ------------- */

table.em-calendar thead { background: #203864; }
table.em-calendar td.eventful-today a , table.em-calendar td.eventful a { color: #203864; }

#tribe-events-content .tribe-events-tooltip h4, #tribe_events_filters_wrapper .tribe_events_slider_val, .single-tribe_events a.tribe-events-ical,
.single-tribe_events a.tribe-events-gcal {
  color: #203864;
  }
.tribe-events-calendar td.tribe-events-present div[id*="tribe-events-daynum-"], .tribe-events-calendar td.tribe-events-present div[id*="tribe-events-daynum-"] > a,
#tribe_events_filters_wrapper input[type=submit], .tribe-events-button, #tribe-events .tribe-events-button, .tribe-events-button.tribe-inactive,
#tribe-events .tribe-events-button:hover, .tribe-events-button:hover, .tribe-events-button.tribe-active:hover {
  background: #203864;
  }

/* ------------ LearnDash LMS --------------*/

#learndash_lessons a, #learndash_quizzes a, .expand_collapse a, .learndash_topic_dots a, .learndash_topic_dots a > span, #learndash_lesson_topics_list span a, #learndash_profile a, #learndash_profile a span {
  color: #203864 !important;
  }
.wpProQuiz_content h2:after { border-color: #203864; }
.wpProQuiz_button, .wpProQuiz_button:hover { background-color: #203864 !important; border-color: #203864 !important; }

/*------- WooCommerce ---------*/

.woocommerce-site .cart-contents .cart-count {
  background: #203864;
}

.woocommerce input[name="update_cart"], .woocommerce input[name="proceed"], .woocommerce input[name="woocommerce_checkout_place_order"],
 .woocommerce-page input[name="update_cart"], .woocommerce-page input[name="proceed"], .woocommerce-page input[name="woocommerce_checkout_place_order"] {
  color: #ffffff;
  background-color: #203864;
  }
.woocommerce a.button, .woocommerce button.button, .woocommerce input.button, .woocommerce #respond input#submit, .woocommerce #content input.button, .woocommerce a.button.alt,
.woocommerce button.button.alt, .woocommerce input.button.alt, .woocommerce #respond input#submit.alt, .woocommerce #content input.button.alt,
.woocommerce-page a.button, .woocommerce-page button.button, .woocommerce-page input.button, .woocommerce-page #respond input#submit,
.woocommerce-page #content input.button, .woocommerce-page a.button.alt, .woocommerce-page button.button.alt, .woocommerce-page input.button.alt,
.woocommerce-page #respond input#submit.alt, .woocommerce-page #content input.button.alt {
background: #203864;
border-color: #203864;
}

.woocommerce a.add_to_cart_button, .woocommerce-page a.add_to_cart_button { background: transparent; border-color: #aaa;}

.woocommerce .quantity .plus, .woocommerce #content .quantity .plus, .woocommerce .quantity .minus, .woocommerce #content .quantity .minus, .woocommerce-page .quantity .plus,
.woocommerce-page #content .quantity .plus, .woocommerce-page .quantity .minus, .woocommerce-page #content .quantity .minus {
background: #203864;
}

.woocommerce .woocommerce-message, .woocommerce .woocommerce-info, .woocommerce .woocommerce-error {
border-color: rgba(32, 56 , 100, 0.3);
background: rgba(32, 56 , 100, 0.1);
}

.woocommerce span.onsale, .woocommerce-page span.onsale { background: #203864; }

.woocommerce-site .cart-contents .cart-count { background: #203864; }

.woocommerce .star-rating span:before, .woocommerce-page .star-rating span:before {
  color: #203864;
  }
.woocommerce span.onsale, .woocommerce-page span.onsale {
  background: #203864;
  text-shadow: none;
  box-shadow: none;
  }
.woocommerce-message,  .woocommerce-info,  .woocommerce-error {
    border: 1px solid rgba(32, 56 , 100, 0.3);
    background: rgba(32, 56 , 100, 0.2);
}
.cart-contents .cart-count {
    background: #203864;
}
ul.products li.product h3:hover {
    color: #203864;
}

.tp_recent_tweets li a { color: #203864 !important; }

.instagram-pics img:hover { border-color: #203864 !important; }

.tp-caption.medium_bg_austin { background-color: #203864 !important; }
.tp-caption.medium_bg_orange { background-color: rgba(32, 56 , 100, 0.75) !important; }

/* =============== END - Skin Styles ============= */

.comments-closed.pings-open {
display: none;
}

.post-snippets .type-post .image-info .terms { display: none; }
</style>
<link rel='stylesheet' id='animate-css-css'  href='http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/animate-css/animate.min.css?ver=5.2' type='text/css' media='all' />
<script type='text/javascript' src='http://www.uees.edu.sv/wp-includes/js/jquery/jquery.js?ver=1.12.4'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-includes/js/jquery/jquery-migrate.min.js?ver=1.4.1'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/easy-video-player/lib/flowplayer.min.js?ver=4.7.5'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/revslider/public/assets/js/jquery.themepunch.tools.min.js?ver=5.4.1'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/revslider/public/assets/js/jquery.themepunch.revolution.min.js?ver=5.4.1'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.easing.1.3.js?ver=4.7.5'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var panelsStyles = {"fullContainer":"body"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/siteorigin-panels/js/styling-263.min.js?ver=2.6.3'></script>
<link rel='https://api.w.org/' href='http://www.uees.edu.sv/?rest_route=/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://www.uees.edu.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://www.uees.edu.sv/wp-includes/wlwmanifest.xml" /> 
<meta name="generator" content="WordPress 4.7.5" />
<link rel='shortlink' href='http://www.uees.edu.sv/' />
<link rel="alternate" type="application/json+oembed" href="http://www.uees.edu.sv/?rest_route=%2Foembed%2F1.0%2Fembed&#038;url=http%3A%2F%2Fwww.uees.edu.sv%2F" />
<link rel="alternate" type="text/xml+oembed" href="http://www.uees.edu.sv/?rest_route=%2Foembed%2F1.0%2Fembed&#038;url=http%3A%2F%2Fwww.uees.edu.sv%2F&#038;format=xml" />
<!-- This content is generated with the Easy Video Player plugin v1.1.7 - http://noorsplugin.com/wordpress-video-plugin/ --><script>flowplayer.conf.embed = false;flowplayer.conf.keyboard = false;</script><!-- Easy Video Player plugin -->            <style type="text/css"></style>            <style type="text/css"></style>            <style type="text/css"></style>            <style type="text/css"></style>            <style type="text/css"></style>            <style type="text/css"></style><meta name="generator" content="Powered by Visual Composer - drag and drop page builder for WordPress."/>
<!--[if lte IE 9]><link rel="stylesheet" type="text/css" href="http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/css/vc_lte_ie9.min.css" media="screen"><![endif]--><meta name="generator" content="Powered by Slider Revolution 5.4.1 - responsive, Mobile-Friendly Slider Plugin for WordPress with comfortable drag and drop interface." />
                <style type="text/css" media="all"
                       id="siteorigin-panels-layouts-head">/* Layout 14611 */ #pgc-14611-0-0 , #pgc-14611-1-0 , #pgc-14611-2-0 , #pgc-14611-3-0 , #pgc-14611-4-0 , #pgc-14611-5-0 , #pgc-14611-6-0 , #pgc-14611-7-0 { width:100%;width:calc(100% - ( 0 * 30px ) ) } #pg-14611-0 , #pg-14611-1 , #pg-14611-2 , #pg-14611-3 , #pg-14611-4 , #pg-14611-5 , #pg-14611-6 , #pg-14611-7 , #pl-14611 .so-panel:last-child { margin-bottom:0px } #pl-14611 .so-panel { margin-bottom:30px } #pg-14611-4> .panel-row-style { background-image:url(http://www.uees.edu.sv/wp-content/uploads/2014/10/geo-bg4.jpg);background-repeat:repeat } #pg-14611-4.panel-no-style, #pg-14611-4.panel-has-style > .panel-row-style { -webkit-align-items:flex-start;align-items:flex-start } #pg-14611-5> .panel-row-style , #pg-14611-6> .panel-row-style { background-color:#eeeeee } @media (max-width:780px){ #pg-14611-0.panel-no-style, #pg-14611-0.panel-has-style > .panel-row-style , #pg-14611-1.panel-no-style, #pg-14611-1.panel-has-style > .panel-row-style , #pg-14611-2.panel-no-style, #pg-14611-2.panel-has-style > .panel-row-style , #pg-14611-3.panel-no-style, #pg-14611-3.panel-has-style > .panel-row-style , #pg-14611-4.panel-no-style, #pg-14611-4.panel-has-style > .panel-row-style , #pg-14611-5.panel-no-style, #pg-14611-5.panel-has-style > .panel-row-style , #pg-14611-6.panel-no-style, #pg-14611-6.panel-has-style > .panel-row-style , #pg-14611-7.panel-no-style, #pg-14611-7.panel-has-style > .panel-row-style { -webkit-flex-direction:column;-ms-flex-direction:column;flex-direction:column } #pg-14611-0 .panel-grid-cell , #pg-14611-1 .panel-grid-cell , #pg-14611-2 .panel-grid-cell , #pg-14611-3 .panel-grid-cell , #pg-14611-4 .panel-grid-cell , #pg-14611-5 .panel-grid-cell , #pg-14611-6 .panel-grid-cell , #pg-14611-7 .panel-grid-cell { margin-right:0 } #pg-14611-0 .panel-grid-cell , #pg-14611-1 .panel-grid-cell , #pg-14611-2 .panel-grid-cell , #pg-14611-3 .panel-grid-cell , #pg-14611-4 .panel-grid-cell , #pg-14611-5 .panel-grid-cell , #pg-14611-6 .panel-grid-cell , #pg-14611-7 .panel-grid-cell { width:100% } #pl-14611 .panel-grid-cell { padding:0 } #pl-14611 .panel-grid .panel-grid-cell-empty { display:none } #pl-14611 .panel-grid .panel-grid-cell-mobile-last { margin-bottom:0px }  } </style><link rel="icon" href="http://www.uees.edu.sv/wp-content/uploads/2017/06/cropped-top-32x32.png" sizes="32x32" />
<link rel="icon" href="http://www.uees.edu.sv/wp-content/uploads/2017/06/cropped-top-192x192.png" sizes="192x192" />
<link rel="apple-touch-icon-precomposed" href="http://www.uees.edu.sv/wp-content/uploads/2017/06/cropped-top-180x180.png" />
<meta name="msapplication-TileImage" content="http://www.uees.edu.sv/wp-content/uploads/2017/06/cropped-top-270x270.png" />

<!-- BEGIN GADWP v5.3.1.1 Universal Analytics - https://deconf.com/google-analytics-dashboard-wordpress/ -->
<script>
(function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
	(i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
	m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
})(window,document,'script','https://www.google-analytics.com/analytics.js','ga');
  ga('create', 'UA-107318580-2', 'auto');
  ga('send', 'pageview');
</script>
<!-- END GADWP Universal Analytics -->
<noscript><style type="text/css"> .wpb_animate_when_almost_visible { opacity: 1; }</style></noscript><style type="text/css">/** Mega Menu CSS: fs **/</style>

</head>

<body class="home page-template page-template-template-1c page-template-template-1c-php page page-id-14611 siteorigin-panels siteorigin-panels-before-js siteorigin-panels-home mega-menu-primary layout-1c  wpb-js-composer js-comp-ver-5.2 vc_responsive">

<div id="page-loading"></div>

<a id="mobile-menu-toggle" href="#"><i class="icon-reorder"></i>&nbsp;</a>
<nav id="mobile-menu" class="menu-container clearfix"><div class="menu-header">Menu</div><div id="mega-menu-wrap-primary" class="mega-menu-wrap"><div class="mega-menu-toggle" tabindex="0"><div class="mega-toggle-blocks-left"><div class='mega-toggle-block mega-menu-toggle-block mega-toggle-block-1' id='mega-toggle-block-1'><span class='mega-toggle-label'><span class='mega-toggle-label-closed'>MENU</span><span class='mega-toggle-label-open'>MENU</span></span></div></div><div class="mega-toggle-blocks-center"></div><div class="mega-toggle-blocks-right"></div></div><ul id="mega-menu-primary" class="mega-menu mega-menu-horizontal mega-no-js" data-event="hover_intent" data-effect="fade" data-effect-speed="200" data-effect-mobile="disabled" data-effect-speed-mobile="200" data-second-click="close" data-document-click="collapse" data-vertical-behaviour="standard" data-breakpoint="800" data-unbind="true"><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-home mega-current-menu-item mega-page_item mega-page-item-14611 mega-current_page_item mega-align-bottom-left mega-menu-flyout mega-item-align-float-left mega-menu-item-15029' id='mega-menu-item-15029'><a class="mega-menu-link" href="http://www.uees.edu.sv/" tabindex="0">Inicio</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-item-align-float-left mega-menu-item-15043' id='mega-menu-item-15043'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=25" aria-haspopup="true" tabindex="0">La Universidad</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-hide-sub-menu-on-mobile mega-menu-item-13778' id='mega-menu-item-13778'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=25">Historia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-hide-sub-menu-on-mobile mega-menu-item-17560' id='mega-menu-item-17560'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17559" aria-haspopup="true">Docencia</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13808' id='mega-menu-item-13808'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=53">Mensaje de Vicerectora Académica</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13792' id='mega-menu-item-13792'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=69">Dirección de Educación Virtual</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13794' id='mega-menu-item-13794'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=67">Planeamiento y Evaluación Curricular</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13804' id='mega-menu-item-13804'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=57">Evaluación y Acreditación</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-17425' id='mega-menu-item-17425'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17424" aria-haspopup="true">Investigación, Proyección Social y Difusión Científica</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13806' id='mega-menu-item-13806'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=55">Mensaje de Vicerrector de Investigación y Proyección Social</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18295' id='mega-menu-item-18295'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18294">Arte y Cultura</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18291' id='mega-menu-item-18291'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18290">Deportes</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17403' id='mega-menu-item-17403'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=326">Proyección Social y Servicios Estudiantiles</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19313' id='mega-menu-item-19313'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17683">Dirección de Publicaciones</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19581' id='mega-menu-item-19581'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19580">Comité de Ética para la Investigación en Salud(CEIS UEES)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17404' id='mega-menu-item-17404'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16411">Dirección de investigación</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13798' id='mega-menu-item-13798'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=63">Organización Institucional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18437' id='mega-menu-item-18437'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18304">Relaciones y Cooperación Internacional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19993' id='mega-menu-item-19993'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19966">Sistema de Gestión de Calidad</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13790' id='mega-menu-item-13790'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=71">Memoria de Labores</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-menu-item-18569' id='mega-menu-item-18569'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279" aria-haspopup="true" tabindex="0">Nuevo Ingreso</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-14231' id='mega-menu-item-14231'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279" aria-haspopup="true">Admisión</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16326' id='mega-menu-item-16326'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279">Matricula</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16175' id='mega-menu-item-16175'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16174">Aranceles</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16328' id='mega-menu-item-16328'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16327">Tramites</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16338' id='mega-menu-item-16338'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16337">Requisitos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16344' id='mega-menu-item-16344'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16343">Calendario Académico</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16354' id='mega-menu-item-16354'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16353">Documentos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16380' id='mega-menu-item-16380'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16379">Admisión a Extranjeros</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15104' id='mega-menu-item-15104'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15103">¿Preguntas frecuentes?</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-19287' id='mega-menu-item-19287'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19260" aria-haspopup="true">Pregrado</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-19261' id='mega-menu-item-19261'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19260" aria-haspopup="true">Facultades</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15567' id='mega-menu-item-15567'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15566" aria-haspopup="true">Facultad de Medicina</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15460' id='mega-menu-item-15460'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15459">Doctorado en Medicina</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15519' id='mega-menu-item-15519'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15518">Licenciatura en Enfermería</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15533' id='mega-menu-item-15533'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15532">Licenciatura  en Nutrición y Dietética</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15547' id='mega-menu-item-15547'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15546">Técnico en Enfermería</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15590' id='mega-menu-item-15590'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15588" aria-haspopup="true">Facultad de Odontología</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15598' id='mega-menu-item-15598'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15596">Doctorado en Cirugía Dental</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15607' id='mega-menu-item-15607'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15606">Técnico en Asistencia Dental</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15695' id='mega-menu-item-15695'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15691" aria-haspopup="true">Facultad de Ingenierías</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15665' id='mega-menu-item-15665'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15664">Ingeniería en Sistemas Computacionales</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15682' id='mega-menu-item-15682'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15680">Técnico en Redes y Tecnologías Informáticas</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15711' id='mega-menu-item-15711'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15709" aria-haspopup="true">Facultad de Ciencias Jurídicas</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15719' id='mega-menu-item-15719'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15718">Licenciatura en Ciencias Jurídicas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15729' id='mega-menu-item-15729'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15724">Licenciatura  en Relaciones y Negocios  Internacionales</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15770' id='mega-menu-item-15770'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15758" aria-haspopup="true">Facultad de Ciencias Sociales</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15784' id='mega-menu-item-15784'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15783">Licenciatura en traducción e Interpretación del Idioma Inglés</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15790' id='mega-menu-item-15790'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15789">Licenciatura en Educación Especial</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15800' id='mega-menu-item-15800'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15798">Licenciatura en Psicología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15809' id='mega-menu-item-15809'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15808">Licenciatura en Teología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15820' id='mega-menu-item-15820'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15819">Licenciatura y Profesorado en educación Parvularia</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15894' id='mega-menu-item-15894'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15892" aria-haspopup="true">Facultad de Ciencias Empresariales y Económicas</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15908' id='mega-menu-item-15908'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15907">Licenciatura en Administración de Empresas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15913' id='mega-menu-item-15913'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15912">Licenciatura en Mercadotecnia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15916' id='mega-menu-item-15916'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15915">Licenciatura en Contaduría Pública</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15922' id='mega-menu-item-15922'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15921">Lic. en Relaciones Públicas con especialidad en Marketing</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15925' id='mega-menu-item-15925'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15924">Técnico en Mercadotecnia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15928' id='mega-menu-item-15928'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15927">Técnico en Relaciones Públicas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15931' id='mega-menu-item-15931'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15930">Técnico/a en Marketing Turístico</a></li>			</ul>
</li>		</ul>
</li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16152' id='mega-menu-item-16152'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16151" aria-haspopup="true">Posgrado UEES</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16300' id='mega-menu-item-16300'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16151" aria-haspopup="true">Maestrías</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21391' id='mega-menu-item-21391'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21390">Posgrado en Gerencia en Salud (Modalidad Semipresencial)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21383' id='mega-menu-item-21383'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21382">Programa de Certificación en Inbound Marketing</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20334' id='mega-menu-item-20334'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20314">Maestría en Epidemiología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16136' id='mega-menu-item-16136'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16135">Maestría en Salud Familiar</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16096' id='mega-menu-item-16096'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16095">Maestría en Derecho de Familia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16155' id='mega-menu-item-16155'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16154">Maestría en Salud Pública</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16141' id='mega-menu-item-16141'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16140">Maestría en Recursos Humanos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16149' id='mega-menu-item-16149'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16147">Maestría en Metodología de la Investigación Cietífica</a></li>		</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-21366' id='mega-menu-item-21366'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21361" aria-haspopup="true">Cursos</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21365' id='mega-menu-item-21365'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21361">Derecho Medioambiental</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21373' id='mega-menu-item-21373'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21372">Curso de Electrocardiografía</a></li>		</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16210' id='mega-menu-item-16210'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16209" aria-haspopup="true">Diplomados</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16239' id='mega-menu-item-16239'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16237" aria-haspopup="true">EPOUEES</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16282' id='mega-menu-item-16282'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16281">Operatoria y Rehabilitacición Oral Avanzada</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16286' id='mega-menu-item-16286'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16285">Odontologia Infantil y Aparatología Interceptiva</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16289' id='mega-menu-item-16289'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16288">Endodoncia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20832' id='mega-menu-item-20832'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20831">Curso de Oclusión aplicada a la Clínica</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20837' id='mega-menu-item-20837'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20836">Implantología y Rehabilitación Bucal</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21388' id='mega-menu-item-21388'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21387">Investigación Científica (Modalidad Virtual)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21380' id='mega-menu-item-21380'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21379">Diplomado en Epidemiología (Modalidad Virtual)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16217' id='mega-menu-item-16217'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16214">Diplomado en Gestión Estratégica del Marketing Digital</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16221' id='mega-menu-item-16221'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16215">Proyecto con enfoque en Salud</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16225' id='mega-menu-item-16225'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16224">Investigación Social</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16231' id='mega-menu-item-16231'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16230">Posgrado de Gerencia en Salud, Semipresencial</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16235' id='mega-menu-item-16235'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16234">Docencia de la Educación Superior (Modalidad Virtual)</a></li>		</ul>
</li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13827' id='mega-menu-item-13827'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=123">Becas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17529' id='mega-menu-item-17529'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17528">Beneficios UEES</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13829' id='mega-menu-item-13829'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=120">Orientación Vocacional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17531' id='mega-menu-item-17531'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=61">Convenios</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-custom mega-menu-item-object-custom mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-menu-item-15871' id='mega-menu-item-15871'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15566" aria-haspopup="true" tabindex="0">Estudiantes</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21522' id='mega-menu-item-21522'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21520">Unidad de Egresados</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15990' id='mega-menu-item-15990'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15989">Portal del Estudiante</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19174' id='mega-menu-item-19174'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19173">Secretaria de Asuntos Espirituales</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13825' id='mega-menu-item-13825'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=126">Reglamentos</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-18109' id='mega-menu-item-18109'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=322" tabindex="0">Portal del Docente</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-20247' id='mega-menu-item-20247'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16448" tabindex="0">Graduados</a></li><li class='mega-menu-item mega-menu-item-type-custom mega-menu-item-object-custom mega-align-bottom-left mega-menu-flyout mega-menu-item-20248' id='mega-menu-item-20248'><a class="mega-menu-link" href="http://ojs.uees.edu.sv/ModU/biblioteca/index2.php" tabindex="0">Biblioteca</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-19393' id='mega-menu-item-19393'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19392" tabindex="0">UEES Virtual</a></li></ul></div></nav><!-- #mobile-menu -->
<div id="container">

    
    
    <header id="header" >

        
        <div class="inner clearfix">

            <div class="wrap">

                <h1 id="site-logo"><a href="http://www.uees.edu.sv/" title="Universidad Evangélica de El Salvador" rel="home"><img class="standard-logo" src="http://www.uees.edu.sv/wp-content/uploads/2017/06/logo140.png" alt="Universidad Evangélica de El Salvador"/></a></h1><nav id="primary-menu" class="dropdown-menu-wrap clearfix"><div id="mega-menu-wrap-primary" class="mega-menu-wrap"><div class="mega-menu-toggle" tabindex="0"><div class="mega-toggle-blocks-left"><div class='mega-toggle-block mega-menu-toggle-block mega-toggle-block-1' id='mega-toggle-block-1'><span class='mega-toggle-label'><span class='mega-toggle-label-closed'>MENU</span><span class='mega-toggle-label-open'>MENU</span></span></div></div><div class="mega-toggle-blocks-center"></div><div class="mega-toggle-blocks-right"></div></div><ul id="mega-menu-primary" class="mega-menu mega-menu-horizontal mega-no-js" data-event="hover_intent" data-effect="fade" data-effect-speed="200" data-effect-mobile="disabled" data-effect-speed-mobile="200" data-second-click="close" data-document-click="collapse" data-vertical-behaviour="standard" data-breakpoint="800" data-unbind="true"><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-home mega-current-menu-item mega-page_item mega-page-item-14611 mega-current_page_item mega-align-bottom-left mega-menu-flyout mega-item-align-float-left mega-menu-item-15029' id='mega-menu-item-15029'><a class="mega-menu-link" href="http://www.uees.edu.sv/" tabindex="0">Inicio</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-item-align-float-left mega-menu-item-15043' id='mega-menu-item-15043'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=25" aria-haspopup="true" tabindex="0">La Universidad</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-hide-sub-menu-on-mobile mega-menu-item-13778' id='mega-menu-item-13778'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=25">Historia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-hide-sub-menu-on-mobile mega-menu-item-17560' id='mega-menu-item-17560'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17559" aria-haspopup="true">Docencia</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13808' id='mega-menu-item-13808'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=53">Mensaje de Vicerectora Académica</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13792' id='mega-menu-item-13792'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=69">Dirección de Educación Virtual</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13794' id='mega-menu-item-13794'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=67">Planeamiento y Evaluación Curricular</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13804' id='mega-menu-item-13804'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=57">Evaluación y Acreditación</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-17425' id='mega-menu-item-17425'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17424" aria-haspopup="true">Investigación, Proyección Social y Difusión Científica</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13806' id='mega-menu-item-13806'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=55">Mensaje de Vicerrector de Investigación y Proyección Social</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18295' id='mega-menu-item-18295'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18294">Arte y Cultura</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18291' id='mega-menu-item-18291'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18290">Deportes</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17403' id='mega-menu-item-17403'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=326">Proyección Social y Servicios Estudiantiles</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19313' id='mega-menu-item-19313'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17683">Dirección de Publicaciones</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19581' id='mega-menu-item-19581'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19580">Comité de Ética para la Investigación en Salud(CEIS UEES)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17404' id='mega-menu-item-17404'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16411">Dirección de investigación</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13798' id='mega-menu-item-13798'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=63">Organización Institucional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-18437' id='mega-menu-item-18437'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=18304">Relaciones y Cooperación Internacional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19993' id='mega-menu-item-19993'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19966">Sistema de Gestión de Calidad</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13790' id='mega-menu-item-13790'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=71">Memoria de Labores</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-menu-item-18569' id='mega-menu-item-18569'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279" aria-haspopup="true" tabindex="0">Nuevo Ingreso</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-14231' id='mega-menu-item-14231'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279" aria-haspopup="true">Admisión</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16326' id='mega-menu-item-16326'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=279">Matricula</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16175' id='mega-menu-item-16175'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16174">Aranceles</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16328' id='mega-menu-item-16328'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16327">Tramites</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16338' id='mega-menu-item-16338'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16337">Requisitos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16344' id='mega-menu-item-16344'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16343">Calendario Académico</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16354' id='mega-menu-item-16354'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16353">Documentos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16380' id='mega-menu-item-16380'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16379">Admisión a Extranjeros</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15104' id='mega-menu-item-15104'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15103">¿Preguntas frecuentes?</a></li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-19287' id='mega-menu-item-19287'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19260" aria-haspopup="true">Pregrado</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-19261' id='mega-menu-item-19261'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19260" aria-haspopup="true">Facultades</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15567' id='mega-menu-item-15567'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15566" aria-haspopup="true">Facultad de Medicina</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15460' id='mega-menu-item-15460'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15459">Doctorado en Medicina</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15519' id='mega-menu-item-15519'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15518">Licenciatura en Enfermería</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15533' id='mega-menu-item-15533'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15532">Licenciatura  en Nutrición y Dietética</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15547' id='mega-menu-item-15547'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15546">Técnico en Enfermería</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15590' id='mega-menu-item-15590'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15588" aria-haspopup="true">Facultad de Odontología</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15598' id='mega-menu-item-15598'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15596">Doctorado en Cirugía Dental</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15607' id='mega-menu-item-15607'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15606">Técnico en Asistencia Dental</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15695' id='mega-menu-item-15695'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15691" aria-haspopup="true">Facultad de Ingenierías</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15665' id='mega-menu-item-15665'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15664">Ingeniería en Sistemas Computacionales</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15682' id='mega-menu-item-15682'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15680">Técnico en Redes y Tecnologías Informáticas</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15711' id='mega-menu-item-15711'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15709" aria-haspopup="true">Facultad de Ciencias Jurídicas</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15719' id='mega-menu-item-15719'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15718">Licenciatura en Ciencias Jurídicas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15729' id='mega-menu-item-15729'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15724">Licenciatura  en Relaciones y Negocios  Internacionales</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15770' id='mega-menu-item-15770'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15758" aria-haspopup="true">Facultad de Ciencias Sociales</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15784' id='mega-menu-item-15784'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15783">Licenciatura en traducción e Interpretación del Idioma Inglés</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15790' id='mega-menu-item-15790'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15789">Licenciatura en Educación Especial</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15800' id='mega-menu-item-15800'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15798">Licenciatura en Psicología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15809' id='mega-menu-item-15809'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15808">Licenciatura en Teología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15820' id='mega-menu-item-15820'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15819">Licenciatura y Profesorado en educación Parvularia</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-15894' id='mega-menu-item-15894'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15892" aria-haspopup="true">Facultad de Ciencias Empresariales y Económicas</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15908' id='mega-menu-item-15908'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15907">Licenciatura en Administración de Empresas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15913' id='mega-menu-item-15913'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15912">Licenciatura en Mercadotecnia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15916' id='mega-menu-item-15916'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15915">Licenciatura en Contaduría Pública</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15922' id='mega-menu-item-15922'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15921">Lic. en Relaciones Públicas con especialidad en Marketing</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15925' id='mega-menu-item-15925'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15924">Técnico en Mercadotecnia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15928' id='mega-menu-item-15928'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15927">Técnico en Relaciones Públicas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15931' id='mega-menu-item-15931'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15930">Técnico/a en Marketing Turístico</a></li>			</ul>
</li>		</ul>
</li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16152' id='mega-menu-item-16152'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16151" aria-haspopup="true">Posgrado UEES</a>
	<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16300' id='mega-menu-item-16300'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16151" aria-haspopup="true">Maestrías</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21391' id='mega-menu-item-21391'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21390">Posgrado en Gerencia en Salud (Modalidad Semipresencial)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21383' id='mega-menu-item-21383'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21382">Programa de Certificación en Inbound Marketing</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20334' id='mega-menu-item-20334'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20314">Maestría en Epidemiología</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16136' id='mega-menu-item-16136'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16135">Maestría en Salud Familiar</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16096' id='mega-menu-item-16096'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16095">Maestría en Derecho de Familia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16155' id='mega-menu-item-16155'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16154">Maestría en Salud Pública</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16141' id='mega-menu-item-16141'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16140">Maestría en Recursos Humanos</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16149' id='mega-menu-item-16149'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16147">Maestría en Metodología de la Investigación Cietífica</a></li>		</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-21366' id='mega-menu-item-21366'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21361" aria-haspopup="true">Cursos</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21365' id='mega-menu-item-21365'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21361">Derecho Medioambiental</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21373' id='mega-menu-item-21373'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21372">Curso de Electrocardiografía</a></li>		</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16210' id='mega-menu-item-16210'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16209" aria-haspopup="true">Diplomados</a>
		<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-has-children mega-menu-item-16239' id='mega-menu-item-16239'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16237" aria-haspopup="true">EPOUEES</a>
			<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16282' id='mega-menu-item-16282'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16281">Operatoria y Rehabilitacición Oral Avanzada</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16286' id='mega-menu-item-16286'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16285">Odontologia Infantil y Aparatología Interceptiva</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16289' id='mega-menu-item-16289'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16288">Endodoncia</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20832' id='mega-menu-item-20832'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20831">Curso de Oclusión aplicada a la Clínica</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-20837' id='mega-menu-item-20837'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=20836">Implantología y Rehabilitación Bucal</a></li>			</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21388' id='mega-menu-item-21388'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21387">Investigación Científica (Modalidad Virtual)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21380' id='mega-menu-item-21380'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21379">Diplomado en Epidemiología (Modalidad Virtual)</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16217' id='mega-menu-item-16217'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16214">Diplomado en Gestión Estratégica del Marketing Digital</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16221' id='mega-menu-item-16221'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16215">Proyecto con enfoque en Salud</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16225' id='mega-menu-item-16225'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16224">Investigación Social</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16231' id='mega-menu-item-16231'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16230">Posgrado de Gerencia en Salud, Semipresencial</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-16235' id='mega-menu-item-16235'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16234">Docencia de la Educación Superior (Modalidad Virtual)</a></li>		</ul>
</li>	</ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13827' id='mega-menu-item-13827'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=123">Becas</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17529' id='mega-menu-item-17529'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=17528">Beneficios UEES</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13829' id='mega-menu-item-13829'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=120">Orientación Vocacional</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-17531' id='mega-menu-item-17531'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=61">Convenios</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-custom mega-menu-item-object-custom mega-menu-item-has-children mega-align-bottom-left mega-menu-flyout mega-menu-item-15871' id='mega-menu-item-15871'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15566" aria-haspopup="true" tabindex="0">Estudiantes</a>
<ul class="mega-sub-menu">
<li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-21522' id='mega-menu-item-21522'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=21520">Unidad de Egresados</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-15990' id='mega-menu-item-15990'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=15989">Portal del Estudiante</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-19174' id='mega-menu-item-19174'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19173">Secretaria de Asuntos Espirituales</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-menu-item-13825' id='mega-menu-item-13825'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=126">Reglamentos</a></li></ul>
</li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-18109' id='mega-menu-item-18109'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=322" tabindex="0">Portal del Docente</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-20247' id='mega-menu-item-20247'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=16448" tabindex="0">Graduados</a></li><li class='mega-menu-item mega-menu-item-type-custom mega-menu-item-object-custom mega-align-bottom-left mega-menu-flyout mega-menu-item-20248' id='mega-menu-item-20248'><a class="mega-menu-link" href="http://ojs.uees.edu.sv/ModU/biblioteca/index2.php" tabindex="0">Biblioteca</a></li><li class='mega-menu-item mega-menu-item-type-post_type mega-menu-item-object-page mega-align-bottom-left mega-menu-flyout mega-menu-item-19393' id='mega-menu-item-19393'><a class="mega-menu-link" href="http://www.uees.edu.sv/?page_id=19392" tabindex="0">UEES Virtual</a></li></ul></div></nav><!-- #primary-menu -->
                
            </div>

        </div>

    </header>
    <!-- #header -->

    
    <div id="slider-area" class="clearfix"><link href="http://fonts.googleapis.com/css?family=Montserrat:700%2C400|Open+Sans:400|Roboto:700" rel="stylesheet" property="stylesheet" type="text/css" media="all">
<div id="rev_slider_25_1_wrapper" class="rev_slider_wrapper fullwidthbanner-container" data-source="gallery" style="margin:0px auto;background:#eeeeee;padding:0px;margin-top:0px;margin-bottom:0px;">
<!-- START REVOLUTION SLIDER 5.4.1 auto mode -->
	<div id="rev_slider_25_1" class="rev_slider fullwidthabanner" style="display:none;" data-version="5.4.1">
<ul>	<!-- SLIDE  -->
	<li data-index="rs-130" data-transition="fade" data-slotamount="7" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="500"  data-thumb="http://localhost/yolia/wp-content/uploads/2015/05/homeslider_thumb1.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Intro" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png"  alt="" title="transparente1"  width="498" height="319" data-lazyload="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/transparent.png" data-bgposition="center top" data-bgfit="cover" data-bgrepeat="no-repeat" data-bgparallax="1" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<a class="tp-caption   tp-resizeme" 
 href="http://www.uees.edu.sv/?page_id=16151" target="_self"			 id="slide-130-layer-1" 
			 data-x="-187" 
			 data-y="9" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":420,"speed":400,"frame":"0","from":"opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":300,"frame":"999","to":"opacity:0;","ease":"Power3.easeInOut"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 5;text-decoration: none;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="1450px" data-hh="658px" width="1024" height="464" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/2017/06/descuentograd_portada1.jpg" data-no-retina> </a>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-73" data-transition="fade" data-slotamount="7" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="500"  data-thumb="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/slidebg1-100x50.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Intro" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png"  alt="" title="Inicio"  data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/slidebg1.jpg" data-bgposition="center top" data-bgfit="cover" data-bgrepeat="no-repeat" data-bgparallax="1" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 2 -->
		<a class="tp-caption   tp-resizeme rs-parallaxlevel-1" 
 href="http://www.uees.edu.sv/?page_id=20268" target="_self"			 id="slide-73-layer-2" 
			 data-x="501" 
			 data-y="63" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":1400,"speed":710,"frame":"0","from":"y:top;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0.75;sY:0.75;skX:0;skY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 5;text-decoration: none;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="auto" data-hh="auto" width="600" height="429" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/2018/01/congreso.png" data-no-retina> </a>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-73-layer-4" 
			 data-x="207" 
			 data-y="143" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2150,"speed":510,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 6; white-space: nowrap; font-size: 50px; font-weight: 700; color: #1f1f1f; letter-spacing: px;">AL </div>

		<!-- LAYER NR. 4 -->
		<div class="tp-caption blackthin342   tp-resizeme" 
			 id="slide-73-layer-6" 
			 data-x="125" 
			 data-y="209" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2350,"speed":500,"frame":"0","from":"x:0;y:100;z:0;rX:0;rY:0;rZ:0;sX:1;sY:3;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Back.easeOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 7; white-space: nowrap; font-size: 40px; font-weight: 700; color: #007aff; letter-spacing: px;">CONGRESO </div>

		<!-- LAYER NR. 5 -->
		<div class="tp-caption   tp-resizeme" 
			 id="slide-73-layer-7" 
			 data-x="33" 
			 data-y="425" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2500,"speed":300,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 8;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="auto" data-hh="auto" width="440" height="2" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/greyline.png" data-no-retina> </div>

		<!-- LAYER NR. 6 -->
		<a class="tp-caption   tp-resizeme" 
 href="http://www.uees.edu.sv/?page_id=20268" target="_self"			 id="slide-73-layer-8" 
			 data-x="148" 
			 data-y="468" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":2900,"speed":510,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 9; white-space: nowrap; font-size: 20px; line-height: 22px; font-weight: 400; color: #ffffff; letter-spacing: 0px;font-family:Open Sans;text-decoration: none;"><button class="btn btn-warning btn-icon-right btn-block btn-lg btn-effect-icon-slide-in" type="button" style="min-height: 0px; min-width: 0px; line-height: 16px; border-width: 1px; margin: 0px; padding: 15px 40px; letter-spacing: 0px; font-size: 15px;"><span style="min-height: 0px; min-width: 0px; line-height: 13px; border-width: 0px; margin: 0px; padding: 0px; letter-spacing: 0px; font-size: 15px;">VER INFOMACIÓN</span></button> </a>

		<!-- LAYER NR. 7 -->
		<div class="tp-caption blackthin342   tp-resizeme" 
			 id="slide-73-layer-9" 
			 data-x="71" 
			 data-y="268" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2350,"speed":500,"frame":"0","from":"x:0;y:100;z:0;rX:0;rY:0;rZ:0;sX:1;sY:3;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Back.easeOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 10; white-space: nowrap; font-size: 40px; font-weight: 700; color: #007aff; letter-spacing: px;"> INTERNACIONAL </div>

		<!-- LAYER NR. 8 -->
		<div class="tp-caption blackthin342   tp-resizeme" 
			 id="slide-73-layer-10" 
			 data-x="178" 
			 data-y="351" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2350,"speed":500,"frame":"0","from":"x:0;y:100;z:0;rX:0;rY:0;rZ:0;sX:1;sY:3;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Back.easeOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 11; white-space: nowrap; font-size: 60px; font-weight: 700; color: #ec971f; letter-spacing: px;">2018 </div>

		<!-- LAYER NR. 9 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-73-layer-11" 
			 data-x="65" 
			 data-y="68" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2150,"speed":510,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 12; white-space: nowrap; font-size: 50px; font-weight: 700; color: #1f1f1f; letter-spacing: px;">BIENVENIDOS </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-137" data-transition="fade" data-slotamount="7" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="500"  data-thumb="http://localhost/yolia/wp-content/uploads/2015/05/homeslider_thumb1.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Intro" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png"  alt="" title="transparente1"  width="498" height="319" data-lazyload="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/transparent.png" data-bgposition="center top" data-bgfit="cover" data-bgrepeat="no-repeat" data-bgparallax="1" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 10 -->
		<a class="tp-caption   tp-resizeme" 
 href="http://www.uees.edu.sv/?page_id=18304" target="_self"			 id="slide-137-layer-1" 
			 data-x="-217" 
			 data-y="1" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":10,"speed":300,"frame":"0","from":"opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":300,"frame":"999","to":"opacity:0;","ease":"Power3.easeInOut"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 5;text-decoration: none;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="1527px" data-hh="692px" width="1024" height="465" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/2017/06/COMUNICADO-DIRCI_1200x500.jpg" data-no-retina> </a>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-129" data-transition="fade" data-slotamount="7" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="500"  data-thumb="http://localhost/yolia/wp-content/uploads/2015/05/homeslider_thumb1.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Oferta" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png"  alt="" title="posgrado12"  width="1024" height="463" data-lazyload="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/transparent.png" data-bgposition="center top" data-bgfit="cover" data-bgrepeat="no-repeat" data-bgparallax="1" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 11 -->
		<div class="tp-caption   tp-resizeme" 
			 id="slide-129-layer-27" 
			 data-x="-251" 
			 data-y="-18" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":1420,"speed":280,"frame":"0","from":"opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":320,"frame":"999","to":"opacity:0;","ease":"Power3.easeInOut"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 5;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="1605px" data-hh="728px" width="1024" height="463" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/2017/06/posgrado12.jpg" data-no-retina> </div>

		<!-- LAYER NR. 12 -->
		<a class="tp-caption   tp-resizeme" 
 href="http://www.uees.edu.sv/?page_id=16151" target="_self"			 id="slide-129-layer-8" 
			 data-x="101" 
			 data-y="839" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":2900,"speed":480,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 6; white-space: nowrap; font-size: 20px; line-height: 22px; font-weight: 400; color: #ffffff; letter-spacing: 0px;font-family:Open Sans;text-decoration: none;"><button class="btn btn-warning btn-icon-right btn-block btn-lg btn-effect-icon-slide-in" type="button" style="min-height: 0px; min-width: 0px; line-height: 16px; border-width: 1px; margin: 0px; padding: 15px 40px; letter-spacing: 0px; font-size: 15px;"><span style="min-height: 0px; min-width: 0px; line-height: 13px; border-width: 0px; margin: 0px; padding: 0px; letter-spacing: 0px; font-size: 15px;">VER OFERTAS</span></button> </a>

		<!-- LAYER NR. 13 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-129-layer-13" 
			 data-x="-50" 
			 data-y="413" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":40,"speed":2640,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 7; white-space: nowrap; font-size: 30px; font-weight: 700; color: #007aff; letter-spacing: px;">Diplomados </div>

		<!-- LAYER NR. 14 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-129-layer-14" 
			 data-x="-52" 
			 data-y="244" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":100,"speed":2560,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:[100%];","mask":"x:inherit;y:inherit;s:inherit;e:inherit;","ease":"Power3.easeInOut"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 8; white-space: nowrap; font-size: 20px; line-height: 20px; font-weight: 700; color: #444444; letter-spacing: px;">Maestría en Salud Familiar<BR>
Maestría en Salud Pública<BR>
Maestría en Recursos Humanos<BR>
Maestría en Metodología de Investigación Científica<BR>
Maestría en Derecho de Familia<BR> </div>

		<!-- LAYER NR. 15 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-129-layer-15" 
			 data-x="-54" 
			 data-y="478" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":100,"speed":2560,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 9; white-space: nowrap; font-size: 20px; line-height: 20px; font-weight: 700; color: #444444; letter-spacing: px;">Diplomado en Gestión Estratégica del Marketing Digital<BR>
Proyecto con enfoque en Salud<BR>
Investigación Social<BR>
Investigación Científica Modalidad Virtual<BR>
Posgrado de Gerencia en Salud, Semipresencial<BR>
Docencia de la Educación Superior<BR> </div>

		<!-- LAYER NR. 16 -->
		<div class="tp-caption blackmontserrat40   tp-resizeme" 
			 id="slide-129-layer-18" 
			 data-x="-51" 
			 data-y="164" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":100,"speed":2560,"frame":"0","from":"x:0;y:0;z:0;rX:0;rY:0;rZ:0;sX:0;sY:0;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":0,"frame":"999","to":"auto:auto;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 10; white-space: nowrap; font-size: 30px; font-weight: 700; color: #007aff; letter-spacing: px;">Maestrías </div>

		<!-- LAYER NR. 17 -->
		<a class="tp-caption   tp-resizeme" 
 href="http://www.uees.edu.sv/?page_id=16151" target="_self"			 id="slide-129-layer-20" 
			 data-x="304" 
			 data-y="108" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":10,"speed":320,"frame":"0","from":"opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":320,"frame":"999","to":"opacity:0;","ease":"Power3.easeInOut"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 11;text-decoration: none;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="815px" data-hh="518px" width="498" height="319" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/2017/06/transparente1.png" data-no-retina> </a>

		<!-- LAYER NR. 18 -->
		<a class="tp-caption rev-btn " 
 href="http://www.uees.edu.sv/?page_id=16151" target="_self"			 id="slide-129-layer-28" 
			 data-x="122" 
			 data-y="628" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="button" 
			data-actions=''
			data-responsive_offset="on" 
			data-responsive="off"
			data-frames='[{"delay":10,"speed":300,"frame":"0","from":"opacity:0;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":300,"frame":"999","to":"opacity:0;","ease":"Power3.easeInOut"},{"frame":"hover","speed":"0","ease":"Linear.easeNone","to":"o:1;rX:0;rY:0;rZ:0;z:0;","style":"c:rgba(0,0,0,1);bg:rgba(255,255,255,1);bs:solid;bw:0 0 0 0;"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[7,7,7,7]"
			data-paddingright="[20,20,20,20]"
			data-paddingbottom="[7,7,7,7]"
			data-paddingleft="[20,20,20,20]"

			style="z-index: 12; white-space: nowrap; font-size: 12px; line-height: 12px; font-weight: 700; color: #ffcc00; letter-spacing: px;font-family:Roboto;background-color:rgba(0,0,0,0.75);border-color:rgba(0,0,0,1);border-radius:30px 30px 30px 30px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;text-decoration: none;">Ver Información </a>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-74" data-transition="slideup" data-slotamount="7" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="1000"  data-thumb="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dbg-100x50.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Oferta" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png"  alt="" title="Inicio"  data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dbg.jpg" data-bgposition="center top" data-bgfit="cover" data-bgrepeat="no-repeat" data-bgparallax="1" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 19 -->
		<div class="tp-caption   tp-resizeme rs-parallaxlevel-9" 
			 id="slide-74-layer-1" 
			 data-x="212" 
			 data-y="-4" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":1100,"speed":1000,"frame":"0","from":"y:top;","to":"o:1;rZ:33;","ease":"Power3.easeInOut"},{"delay":"+5900","speed":1000,"frame":"999","to":"x:-200px;skX:85px;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 5;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="698px" data-hh="610px" width="800" height="700" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dlayer_6.png" data-no-retina> </div>

		<!-- LAYER NR. 20 -->
		<div class="tp-caption   tp-resizeme rs-parallaxlevel-9" 
			 id="slide-74-layer-2" 
			 data-x="-89" 
			 data-y="-58" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":1400,"speed":1000,"frame":"0","from":"y:top;","to":"o:1;rZ:36;","ease":"Power3.easeInOut"},{"delay":"+5900","speed":1000,"frame":"999","to":"x:-200px;skX:85px;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 6;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="662px" data-hh="539px" width="800" height="700" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dlayer_5.png" data-no-retina> </div>

		<!-- LAYER NR. 21 -->
		<div class="tp-caption   tp-resizeme rs-parallaxlevel-9" 
			 id="slide-74-layer-3" 
			 data-x="-64" 
			 data-y="306" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":1700,"speed":1000,"frame":"0","from":"y:top;","to":"o:1;rZ:32;","ease":"Power3.easeInOut"},{"delay":"+5850","speed":1000,"frame":"999","to":"x:-200px;skX:85px;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 7;"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="637px" data-hh="565px" width="800" height="700" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dlayer_4.png" data-no-retina> </div>

		<!-- LAYER NR. 22 -->
		<div class="tp-caption   tp-resizeme rs-parallaxlevel-3" 
			 id="slide-74-layer-4" 
			 data-x="-256" 
			 data-y="93" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2000,"speed":1000,"frame":"0","from":"y:top;","to":"o:1;rZ:19;","ease":"Power3.easeInOut"},{"delay":"+5900","speed":1000,"frame":"999","to":"x:-200px;skX:85px;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 8;">
<div class="rs-looped rs-slideloop"  data-easing="Linear.easeNone" data-speed="3" data-xs="0" data-xe="0" data-ys="-3" data-ye="3"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="652px" data-hh="575px" width="800" height="700" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dlayer_3.png" data-no-retina> </div></div>

		<!-- LAYER NR. 23 -->
		<div class="tp-caption   tp-resizeme rs-parallaxlevel-1" 
			 id="slide-74-layer-6" 
			 data-x="159" 
			 data-y="220" 
						data-width="['none','none','none','none']"
			data-height="['none','none','none','none']"
 
			data-type="image" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2600,"speed":1000,"frame":"0","from":"y:top;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"+5900","speed":1000,"frame":"999","to":"x:-200px;skX:85px;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 10;">
<div class="rs-looped rs-slideloop"  data-easing="Linear.easeNone" data-speed="2" data-xs="0" data-xe="0" data-ys="-5" data-ye="5"><img src="http://www.uees.edu.sv/wp-content/plugins/revslider/admin/assets/images/dummy.png" alt="" data-ww="613px" data-hh="509px" width="800" height="700" data-lazyload="http://www.uees.edu.sv/wp-content/uploads/revslider/homeslider1/3dlayer_1.png" data-no-retina> </div></div>

		<!-- LAYER NR. 24 -->
		<div class="tp-caption lightmontserrat70shadowed   tp-resizeme rs-parallaxlevel-10" 
			 id="slide-74-layer-7" 
			 data-x="656" 
			 data-y="-6" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2900,"speed":1000,"frame":"0","from":"x:right;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 11; white-space: nowrap; font-size: 50px; color: #ffffff; letter-spacing: px;">CONOCE  </div>

		<!-- LAYER NR. 25 -->
		<div class="tp-caption blackmontserrat60   tp-resizeme rs-parallaxlevel-10" 
			 id="slide-74-layer-8" 
			 data-x="822" 
			 data-y="113" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":3000,"split":"chars","split_direction":"forward","splitdelay":0.1,"speed":1000,"frame":"0","from":"x:0;y:100;z:0;rX:0;rY:0;rZ:0;sX:1;sY:3;skX:0;skY:0;opacity:0;","to":"o:1;","ease":"Power4.easeOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 12; white-space: nowrap; font-weight: 400; color: #1f1f1f; letter-spacing: px;">OFERTA </div>

		<!-- LAYER NR. 26 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15588" target="_self"			 id="slide-74-layer-9" 
			 data-x="808" 
			 data-y="285" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3500,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 13; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE ODONTOLOGÍA </a>

		<!-- LAYER NR. 27 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15691" target="_self"			 id="slide-74-layer-10" 
			 data-x="809" 
			 data-y="335" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3600,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 14; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE INGENIERIAS </a>

		<!-- LAYER NR. 28 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15709" target="_self"			 id="slide-74-layer-11" 
			 data-x="809" 
			 data-y="384" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3700,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 15; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE CIENCIAS JURIDICAS </a>

		<!-- LAYER NR. 29 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15758" target="_self"			 id="slide-74-layer-12" 
			 data-x="808" 
			 data-y="426" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3800,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 16; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE CIENCIAS SOCIALES </a>

		<!-- LAYER NR. 30 -->
		<a class="tp-caption blackboldbgmontserrat207ccedf   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=19260" target="_self"			 id="slide-74-layer-13" 
			 data-x="855" 
			 data-y="530" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3900,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 17; white-space: nowrap; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(124, 206, 223, 1);text-decoration: none;">VER MÁS </a>

		<!-- LAYER NR. 31 -->
		<div class="tp-caption lightmontserrat70shadowed   tp-resizeme rs-parallaxlevel-10" 
			 id="slide-74-layer-15" 
			 data-x="767" 
			 data-y="53" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2900,"speed":1000,"frame":"0","from":"x:right;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 18; white-space: nowrap; font-size: 50px; color: #ffffff; letter-spacing: px;">NUESTRA </div>

		<!-- LAYER NR. 32 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15566" target="_self"			 id="slide-74-layer-16" 
			 data-x="809" 
			 data-y="239" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":8600,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 19; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE MEDICINA </a>

		<!-- LAYER NR. 33 -->
		<a class="tp-caption blackboldbgmontserrat20   tp-resizeme rs-parallaxlevel-10" 
 href="http://www.uees.edu.sv/?page_id=15892" target="_self"			 id="slide-74-layer-17" 
			 data-x="808" 
			 data-y="470" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-actions=''
			data-responsive_offset="on" 

			data-frames='[{"delay":3500,"speed":1000,"frame":"0","from":"x:right;skX:-85px;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[5,5,5,5]"
			data-paddingright="[8,8,8,8]"
			data-paddingbottom="[5,5,5,5]"
			data-paddingleft="[8,8,8,8]"

			style="z-index: 20; white-space: nowrap; font-size: 15px; font-weight: 400; color: #ffffff; letter-spacing: px;background-color:rgba(0, 0, 0, 1);text-decoration: none;">FACULTAD DE CIENCIAS EMPRESARIALES </a>

		<!-- LAYER NR. 34 -->
		<div class="tp-caption lightmontserrat70shadowed   tp-resizeme rs-parallaxlevel-10" 
			 id="slide-74-layer-18" 
			 data-x="726" 
			 data-y="167" 
						data-width="['auto']"
			data-height="['auto']"
 
			data-type="text" 
			data-responsive_offset="on" 

			data-frames='[{"delay":2900,"speed":1000,"frame":"0","from":"x:right;","to":"o:1;","ease":"Power3.easeInOut"},{"delay":"wait","speed":1000,"frame":"999","to":"x:{-250,250};y:{-150,150};rX:{-90,90};rY:{-90,90};rZ:{-360,360};sX:0;sY:0;opacity:0;","ease":"nothing"}]'
			data-textAlign="['inherit','inherit','inherit','inherit']"
			data-paddingtop="[0,0,0,0]"
			data-paddingright="[0,0,0,0]"
			data-paddingbottom="[0,0,0,0]"
			data-paddingleft="[0,0,0,0]"

			style="z-index: 21; white-space: nowrap; font-size: 50px; color: #ffffff; letter-spacing: px;">ACADÉMICA </div>
	</li>
</ul>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss="";
						if(htmlDiv) {
							htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
						}else{
							var htmlDiv = document.createElement("div");
							htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
							document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
						}
					</script>
<div class="tp-bannertimer" style="height: 5px; background: rgba(0,0,0,0.15);"></div>	</div>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss=".tp-caption.blackmontserrat60,.blackmontserrat60{font-size:60px;line-height:60px;font-weight:900;font-family:Montserrat;color:rgb(31,31,31);text-decoration:none;background-color:transparent;border-width:0px;border-color:rgb(0,0,0);border-style:none;text-shadow:none}.tp-caption.blackmontserrat40,.blackmontserrat40{font-size:40px;line-height:40px;font-weight:800;font-family:Montserrat;color:rgb(31,31,31);text-decoration:none;background-color:transparent;border-width:0px;border-color:rgb(31,31,31);border-style:none;text-shadow:none}.tp-caption.blackthin342,.blackthin342{font-size:35px;line-height:35px;font-weight:400;font-family:Montserrat;color:rgb(236,151,31);text-decoration:none;background-color:transparent;border-width:0px;border-color:rgb(0,0,0);border-style:none;text-shadow:none}.tp-caption.lightmontserrat70shadowed,.lightmontserrat70shadowed{font-size:70px;line-height:70px;font-weight:400;font-family:Montserrat;color:rgb(255,255,255);text-decoration:none;background-color:transparent;border-width:0px;border-color:rgb(0,0,0);border-style:none;text-shadow:0px 0px 7px rgba(0,0,0,0.25)}.tp-caption.blackboldbgmontserrat20,.blackboldbgmontserrat20{font-size:20px;line-height:20px;font-weight:900;font-family:Montserrat;color:rgb(255,255,255);text-decoration:none;background-color:rgb(0,0,0);border-width:0px;border-color:rgb(0,0,0);border-style:none;text-shadow:none}.tp-caption.blackboldbgmontserrat207ccedf,.blackboldbgmontserrat207ccedf{font-size:20px;line-height:20px;font-weight:900;font-family:Montserrat;color:rgb(255,255,255);text-decoration:none;background-color:rgb(124,206,223);border-width:0px;border-color:rgb(0,0,0);border-style:none;text-shadow:none}";
				if(htmlDiv) {
					htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
				}else{
					var htmlDiv = document.createElement("div");
					htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
					document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
				}
			</script>
		<script type="text/javascript">
						/******************************************
				-	PREPARE PLACEHOLDER FOR SLIDER	-
			******************************************/

			var setREVStartSize=function(){
				try{var e=new Object,i=jQuery(window).width(),t=9999,r=0,n=0,l=0,f=0,s=0,h=0;
					e.c = jQuery('#rev_slider_25_1');
					e.gridwidth = [1170];
					e.gridheight = [700];
							
					e.sliderLayout = "auto";
					if(e.responsiveLevels&&(jQuery.each(e.responsiveLevels,function(e,f){f>i&&(t=r=f,l=e),i>f&&f>r&&(r=f,n=e)}),t>r&&(l=n)),f=e.gridheight[l]||e.gridheight[0]||e.gridheight,s=e.gridwidth[l]||e.gridwidth[0]||e.gridwidth,h=i/s,h=h>1?1:h,f=Math.round(h*f),"fullscreen"==e.sliderLayout){var u=(e.c.width(),jQuery(window).height());if(void 0!=e.fullScreenOffsetContainer){var c=e.fullScreenOffsetContainer.split(",");if (c) jQuery.each(c,function(e,i){u=jQuery(i).length>0?u-jQuery(i).outerHeight(!0):u}),e.fullScreenOffset.split("%").length>1&&void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0?u-=jQuery(window).height()*parseInt(e.fullScreenOffset,0)/100:void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0&&(u-=parseInt(e.fullScreenOffset,0))}f=u}else void 0!=e.minHeight&&f<e.minHeight&&(f=e.minHeight);e.c.closest(".rev_slider_wrapper").css({height:f})
					
				}catch(d){console.log("Failure at Presize of Slider:"+d)}
			};
			
			setREVStartSize();
			
						var tpj=jQuery;
			tpj.noConflict();
			var revapi25;
			tpj(document).ready(function() {
				if(tpj("#rev_slider_25_1").revolution == undefined){
					revslider_showDoubleJqueryError("#rev_slider_25_1");
				}else{
					revapi25 = tpj("#rev_slider_25_1").show().revolution({
						sliderType:"standard",
jsFileLocation:"//www.uees.edu.sv/wp-content/plugins/revslider/public/assets/js/",
						sliderLayout:"auto",
						dottedOverlay:"none",
						delay:10000,
						navigation: {
							keyboardNavigation:"off",
							keyboard_direction: "horizontal",
							mouseScrollNavigation:"off",
 							mouseScrollReverse:"default",
							onHoverStop:"off",
							touch:{
								touchenabled:"on",
								touchOnDesktop:"off",
								swipe_threshold: 0.7,
								swipe_min_touches: 1,
								swipe_direction: "horizontal",
								drag_block_vertical: false
							}
							,
							arrows: {
								style:"hermes",
								enable:true,
								hide_onmobile:false,
								hide_onleave:false,
								tmp:'<div class="tp-arr-allwrapper">	<div class="tp-arr-imgholder"></div>	<div class="tp-arr-titleholder">{{title}}</div>	</div>',
								left: {
									h_align:"left",
									v_align:"center",
									h_offset:20,
									v_offset:0
								},
								right: {
									h_align:"right",
									v_align:"center",
									h_offset:20,
									v_offset:0
								}
							}
							,
							bullets: {
								enable:true,
								hide_onmobile:false,
								style:"hermes",
								hide_onleave:false,
								direction:"horizontal",
								h_align:"center",
								v_align:"bottom",
								h_offset:0,
								v_offset:20,
								space:5,
								tmp:''
							}
						},
						visibilityLevels:[1240,1024,778,480],
						gridwidth:1170,
						gridheight:700,
						lazyType:"all",
						parallax: {
							type:"mouse",
							origo:"enterpoint",
							speed:400,
							levels:[7,4,3,2,5,4,3,2,1,0,47,48,49,50,51,55],
						},
						shadow:0,
						spinner:"spinner3",
						stopLoop:"off",
						stopAfterLoops:-1,
						stopAtSlide:-1,
						shuffle:"off",
						autoHeight:"off",
						hideThumbsOnMobile:"off",
						hideSliderAtLimit:0,
						hideCaptionAtLimit:0,
						hideAllCaptionAtLilmit:0,
						debugMode:false,
						fallbacks: {
							simplifyAll:"off",
							nextSlideOnWindowFocus:"off",
							disableFocusListener:false,
						}
					});
				}
			});	/*ready*/
		</script>
		<script>
					var htmlDivCss = '	#rev_slider_25_1_wrapper .tp-loader.spinner3 div { background-color: #fff !important; } ';
					var htmlDiv = document.getElementById('rs-plugin-settings-inline-css');
					if(htmlDiv) {
						htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
					}
					else{
						var htmlDiv = document.createElement('div');
						htmlDiv.innerHTML = '<style>' + htmlDivCss + '</style>';
						document.getElementsByTagName('head')[0].appendChild(htmlDiv.childNodes[0]);
					}
					</script>
					<script>
					var htmlDivCss = unescape(".hermes.tparrows%20%7B%0A%09cursor%3Apointer%3B%0A%09background%3Argba%280%2C0%2C0%2C0.5%29%3B%0A%09width%3A30px%3B%0A%09height%3A110px%3B%0A%09position%3Aabsolute%3B%0A%09display%3Ablock%3B%0A%09z-index%3A100%3B%0A%7D%0A%0A.hermes.tparrows%3Abefore%20%7B%0A%09font-family%3A%20%22revicons%22%3B%0A%09font-size%3A15px%3B%0A%09color%3Argb%28255%2C%20255%2C%20255%29%3B%0A%09display%3Ablock%3B%0A%09line-height%3A%20110px%3B%0A%09text-align%3A%20center%3B%0A%20%20%20%20transform%3Atranslatex%280px%29%3B%0A%20%20%20%20-webkit-transform%3Atranslatex%280px%29%3B%0A%20%20%20%20transition%3Aall%200.3s%3B%0A%20%20%20%20-webkit-transition%3Aall%200.3s%3B%0A%7D%0A.hermes.tparrows.tp-leftarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce824%22%3B%0A%7D%0A.hermes.tparrows.tp-rightarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce825%22%3B%0A%7D%0A.hermes.tparrows.tp-leftarrow%3Ahover%3Abefore%20%7B%0A%20%20%20%20transform%3Atranslatex%28-20px%29%3B%0A%20%20%20%20-webkit-transform%3Atranslatex%28-20px%29%3B%0A%20%20%20%20%20opacity%3A0%3B%0A%7D%0A.hermes.tparrows.tp-rightarrow%3Ahover%3Abefore%20%7B%0A%20%20%20%20transform%3Atranslatex%2820px%29%3B%0A%20%20%20%20-webkit-transform%3Atranslatex%2820px%29%3B%0A%20%20%20%20%20opacity%3A0%3B%0A%7D%0A%0A.hermes%20.tp-arr-allwrapper%20%7B%0A%20%20%20%20overflow%3Ahidden%3B%0A%20%20%20%20position%3Aabsolute%3B%0A%09width%3A180px%3B%0A%20%20%20%20height%3A140px%3B%0A%20%20%20%20top%3A0px%3B%0A%20%20%20%20left%3A0px%3B%0A%20%20%20%20visibility%3Ahidden%3B%0A%20%20%20%20%20%20-webkit-transition%3A%20-webkit-transform%200.3s%200.3s%3B%0A%20%20transition%3A%20transform%200.3s%200.3s%3B%0A%20%20-webkit-perspective%3A%201000px%3B%0A%20%20perspective%3A%201000px%3B%0A%20%20%20%20%7D%0A.hermes.tp-rightarrow%20.tp-arr-allwrapper%20%7B%0A%20%20%20right%3A0px%3Bleft%3Aauto%3B%0A%20%20%20%20%20%20%7D%0A.hermes.tparrows%3Ahover%20.tp-arr-allwrapper%20%7B%0A%20%20%20visibility%3Avisible%3B%0A%20%20%20%20%20%20%20%20%20%20%7D%0A.hermes%20.tp-arr-imgholder%20%7B%0A%20%20width%3A180px%3Bposition%3Aabsolute%3B%0A%20%20left%3A0px%3Btop%3A0px%3Bheight%3A110px%3B%0A%20%20transform%3Atranslatex%28-180px%29%3B%0A%20%20-webkit-transform%3Atranslatex%28-180px%29%3B%0A%20%20transition%3Aall%200.3s%3B%0A%20%20transition-delay%3A0.3s%3B%0A%7D%0A.hermes.tp-rightarrow%20.tp-arr-imgholder%7B%0A%20%20%20%20transform%3Atranslatex%28180px%29%3B%0A%20%20-webkit-transform%3Atranslatex%28180px%29%3B%0A%20%20%20%20%20%20%7D%0A%20%20%0A.hermes.tparrows%3Ahover%20.tp-arr-imgholder%20%7B%0A%20%20%20transform%3Atranslatex%280px%29%3B%0A%20%20%20-webkit-transform%3Atranslatex%280px%29%3B%20%20%20%20%20%20%20%20%20%20%20%20%0A%7D%0A.hermes%20.tp-arr-titleholder%20%7B%0A%20%20top%3A110px%3B%0A%20%20width%3A180px%3B%0A%20%20text-align%3Aleft%3B%20%0A%20%20display%3Ablock%3B%0A%20%20padding%3A0px%2010px%3B%0A%20%20line-height%3A30px%3B%20background%3A%23000%3B%0A%20%20background%3Argba%280%2C0%2C0%2C0.75%29%3B%0A%20%20color%3Argb%28255%2C%20255%2C%20255%29%3B%0A%20%20font-weight%3A600%3B%20position%3Aabsolute%3B%0A%20%20font-size%3A12px%3B%0A%20%20white-space%3Anowrap%3B%0A%20%20letter-spacing%3A1px%3B%0A%20%20-webkit-transition%3A%20all%200.3s%3B%0A%20%20transition%3A%20all%200.3s%3B%0A%20%20-webkit-transform%3A%20rotatex%28-90deg%29%3B%0A%20%20transform%3A%20rotatex%28-90deg%29%3B%0A%20%20-webkit-transform-origin%3A%2050%25%200%3B%0A%20%20transform-origin%3A%2050%25%200%3B%0A%20%20box-sizing%3Aborder-box%3B%0A%0A%7D%0A.hermes.tparrows%3Ahover%20.tp-arr-titleholder%20%7B%0A%20%20%20%20-webkit-transition-delay%3A%200.6s%3B%0A%20%20transition-delay%3A%200.6s%3B%0A%20%20-webkit-transform%3A%20rotatex%280deg%29%3B%0A%20%20transform%3A%20rotatex%280deg%29%3B%0A%7D%0A%0A.hermes.tp-bullets%20%7B%0A%7D%0A%0A.hermes%20.tp-bullet%20%7B%0A%20%20%20%20overflow%3Ahidden%3B%0A%20%20%20%20border-radius%3A50%25%3B%0A%20%20%20%20width%3A16px%3B%0A%20%20%20%20height%3A16px%3B%0A%20%20%20%20background-color%3A%20rgba%280%2C%200%2C%200%2C%200%29%3B%0A%20%20%20%20box-shadow%3A%20inset%200%200%200%202px%20rgb%28255%2C%20255%2C%20255%29%3B%0A%20%20%20%20-webkit-transition%3A%20background%200.3s%20ease%3B%0A%20%20%20%20transition%3A%20background%200.3s%20ease%3B%0A%20%20%20%20position%3Aabsolute%3B%0A%7D%0A%0A.hermes%20.tp-bullet%3Ahover%20%7B%0A%09%20%20background-color%3A%20rgba%280%2C0%2C0%2C0.21%29%3B%0A%7D%0A.hermes%20.tp-bullet%3Aafter%20%7B%0A%20%20content%3A%20%27%20%27%3B%0A%20%20position%3A%20absolute%3B%0A%20%20bottom%3A%200%3B%0A%20%20height%3A%200%3B%0A%20%20left%3A%200%3B%0A%20%20width%3A%20100%25%3B%0A%20%20background-color%3A%20rgb%28255%2C%20255%2C%20255%29%3B%0A%20%20box-shadow%3A%200%200%201px%20rgb%28255%2C%20255%2C%20255%29%3B%0A%20%20-webkit-transition%3A%20height%200.3s%20ease%3B%0A%20%20transition%3A%20height%200.3s%20ease%3B%0A%7D%0A.hermes%20.tp-bullet.selected%3Aafter%20%7B%0A%20%20height%3A100%25%3B%0A%7D%0A%0A");
					var htmlDiv = document.getElementById('rs-plugin-settings-inline-css');
					if(htmlDiv) {
						htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
					}
					else{
						var htmlDiv = document.createElement('div');
						htmlDiv.innerHTML = '<style>' + htmlDivCss + '</style>';
						document.getElementsByTagName('head')[0].appendChild(htmlDiv.childNodes[0]);
					}
				  </script>
				</div><!-- END REVOLUTION SLIDER --></div> <!-- #slider-area -->
    <div id="main" class="clearfix">

        
        <div class="inner clearfix">
    <div id="one-column-template" class="layout-1c">

        

    <div id="content" class="twelvecol ">

        
        
            
                
                <article id="post-14611" class="post-14611 page type-page status-publish hentry">

                    
                    <div class="entry-content">

                        
                        <div id="pl-14611"  class="panel-layout" ><div id="pg-14611-0"  class="panel-grid panel-has-style" ><div id="college-intro" class="panel-row-style panel-row-style-for-14611-0" ><div id="pgc-14611-0-0"  class="panel-grid-cell" ><div id="panel-14611-0-0-0" class="so-panel widget widget_mo-heading panel-first-child" data-index="0" ><div class="so-widget-mo-heading so-widget-mo-heading-default-d75171398898">
<div class="heading1 separator"><h3 class="title"><br /><br />Bienvenidos a la Universidad Evangélica de El Salvador</h3></div></div></div><div id="panel-14611-0-0-1" class="so-panel widget widget_mo-tab-slider panel-last-child" data-index="1" ><div class="so-widget-mo-tab-slider so-widget-mo-tab-slider-default-d75171398898"><script type="text/javascript">
jQuery(document).ready(function($) {jQuery('#tab-slider5ab2a4c09f3c9 .flexslider').flexslider({animation: "slide",slideshowSpeed: 5000,animationSpeed: 600,namespace: "flex-",controlNav: true,directionNav: false,smoothHeight: false,animationLoop: false,slideshow: false,easing: "swing",manualControls: "#tab-slider-nav5ab2a4c09f3c9.tab-list li a",controlsContainer: "#tab-slider-nav5ab2a4c09f3c9.tab-list"})});
</script>
<ul id="tab-slider-nav5ab2a4c09f3c9" class="tab-list"><li><a href="#services1">Mensajes</a></li><li><a href="#services2">Catálogo Institucional</a></li><li><a href="#services3">Modelo Educativo</a></li><li><a href="#services4">Convenios</a></li></ul><div id="tab-slider5ab2a4c09f3c9" class="flex-slider-container loading"><div class="flexslider"><ul class="slides"><li id="services1" data-name="Mensajes"><div class="sixcol"><img class="alignnone size-full wp-image-19791" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/FOTOGRAFIARECTOR11.jpg" alt="" width="400" height="300" /></div><div class="sixcol last"><h4>Mensaje de Bienvenida</h4><p>Estimados Estudiantes:</p><p style="text-align: justify;">Las bases filosóficas y pedagógicas de nuestro proyecto educativo nos han orientado desde la fundación de la Universidad en 1981, a asumir los retos y compromisos de la Educación Superior en El Salvador. Esto significa para nosotros el reconocimiento de la importancia fundamental que este tipo de educación reviste para el desarrollo sociocultural y económico de nuestro país y para la construcción del futuro.</p><a class= "button  theme" href="http://www.uees.edu.sv/?page_id=51" target="_self">Ver más</a></div><div class="clear"></div></li><li id="services2" data-name="Catálogo Institucional"><div class="sixcol"><img class="alignnone wp-image-14054" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/bg-contact1.jpg" alt="" width="1108" height="623" /></div><div class="sixcol last"><h4>Catálogo Institucional</h4><p style="text-align: justify;">La Universidad Evangélica de El Salvador (UEES) fue fundada en 1981 por un grupo de cristianos evangélicos, profesionales, líderes de las iglesias evangélicas históricas más representativas de nuestro país (Bautista, Centroamericana y Asambleas de Dios), con un modelo educativo cuyo trasfondo obedece a una cosmovisión bíblica de la historia, el pensamiento y el conocimiento.</p><a class= "button  theme" href="http://www.uees.edu.sv/wp-content/uploads/2017/anunciosFlip/catalogo_institucional/index.html" target="_self">Ver más</a></div><div class="clear"></div></li><li id="services3" data-name="Modelo Educativo"><div class="sixcol"><img class="alignnone wp-image-14057" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/bg-contact3.jpg" alt="" width="1032" height="580" /></div><div class="sixcol last"><h4>Modelo Educativo</h4><p style="text-align: justify;">El Modelo Educativo es un instrumento que contiene las intencionalidades bajo las cuales, la institución, se compromete ante la sociedad en la responsable tarea de formar nuevos cuadros de profesionales en diferentes campos disciplinarios. Su función no sólo orienta la práctica educativa como tarea fundamental, sino las tareas de gestión, administración, desarrollo y evaluación de su quehacer académico y administrativo.</p><a class= "button  theme" href="http://www.uees.edu.sv/wp-content/uploads/2017/anunciosFlip/modelos_educativos/index.html" target="_self">Ver más</a></div><div class="clear"></div></li><li id="services4" data-name="Convenios"><div class="sixcol"><img class="alignnone wp-image-14058" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/bg-contact4.jpg" alt="" width="1039" height="584" /></div><div class="sixcol last"><h4>Convenios</h4><p style="text-align: justify;">La Universidad Evangélica de El Salvador, con el objeto de fortalecer la formación integral y competencia de los miembros de la comunidad educativa, promueve el establecimiento de alianzas estratégicas a nivel nacional, regional e internacional, mediante la suscripción de Convenios y Cartas de Entendimiento.</p><p>.</p><a class= "button  theme" href="http://www.uees.edu.sv/?page_id=61" target="_self">Ver más</a></div><div class="clear"></div></li></ul></div><!-- flexslider --></div><!-- flex-slider-container --></div></div></div></div></div><div id="pg-14611-1"  class="panel-grid panel-has-style" ><div id="college-intro" class="panel-row-style panel-row-style-for-14611-1" ><div id="pgc-14611-1-0"  class="panel-grid-cell" ><div id="panel-14611-1-0-0" class="so-panel widget widget_mo-heading panel-first-child" data-index="2" ><div class="so-widget-mo-heading so-widget-mo-heading-default-d75171398898">
<div class="heading1 separator"><h3 class="title"><br /><br />NOTICIAS Y EVENTOS UEES</h3></div></div></div><div id="panel-14611-1-0-1" class="so-panel widget widget_mo-post-snippets-carousel" data-index="3" ><div class="so-widget-mo-post-snippets-carousel so-widget-mo-post-snippets-carousel-default-d75171398898"><script type="text/javascript">
jQuery(document).ready(function($) {jQuery('#news-carousel .slides').owlCarousel({navigation: false,navigationText: ["<i class=\"icon-uniF489\"></i>","<i class=\"icon-uniF488\"></i>"],scrollPerPage: false,items: 4,itemsDesktop: [1199,4],itemsDesktopSmall: [979,5],itemsTablet: [768,4],itemsTabletSmall: [640,2],itemsMobile: [479,1],autoPlay: 5000,stopOnHover: true,pagination: false,rewindSpeed: 1000,slideSpeed: 200,paginationSpeed: "800"})});
</script>
<div class="carousel-wrap"><div id ="news-carousel" class="carousel-container"><div class="slides image-grid post-snippets  owl-carousel"><article class="post-21472 news type-news status-publish has-post-thumbnail hentry"><div class="image-area"><a title="LA VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL A TRAVÉS DE LA UNIDAD DE ARTE, CULTURA Y DEPORTE, INVITA A PARTICIPAR EN SUS DIFERENTES ACTIVIDADES Y TALLERES" href="http://www.uees.edu.sv/?news=la-vicerrectoria-investigacion-proyeccion-social-traves-la-unidad-arte-cultula-deporte-invita-participar-diferentes-actividades-talleres "><img width="800" height="640" src="http://www.uees.edu.sv/wp-content/uploads/2018/03/AficheTalleres2018.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/03/AficheTalleres2018.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2018/03/AficheTalleres2018-300x240.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2018/03/AficheTalleres2018-768x614.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="LA VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL A TRAVÉS DE LA UNIDAD DE ARTE, CULTURA Y DEPORTE, INVITA A PARTICIPAR EN SUS DIFERENTES ACTIVIDADES Y TALLERES" href="http://www.uees.edu.sv/?news=la-vicerrectoria-investigacion-proyeccion-social-traves-la-unidad-arte-cultula-deporte-invita-participar-diferentes-actividades-talleres ">LA VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL A TRAVÉS DE LA UNIDAD DE ARTE, CULTURA Y DEPORTE, INVITA A PARTICIPAR EN SUS DIFERENTES ACTIVIDADES Y TALLERES</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="LA VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL A TRAVÉS DE LA UNIDAD DE ARTE, CULTURA Y DEPORTE, INVITA A PARTICIPAR EN SUS DIFERENTES ACTIVIDADES Y TALLERES" href="http://www.uees.edu.sv/wp-content/uploads/2018/03/AficheTalleres2018.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=la-vicerrectoria-investigacion-proyeccion-social-traves-la-unidad-arte-cultula-deporte-invita-participar-diferentes-actividades-talleres" title="LA VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL A TRAVÉS DE LA UNIDAD DE ARTE, CULTURA Y DEPORTE, INVITA A PARTICIPAR EN SUS DIFERENTES ACTIVIDADES Y TALLERES">Details</a></div></div></div></article><!-- .hentry --><article class="post-20987 news type-news status-publish has-post-thumbnail hentry"><div class="image-area"><a title="Estudiante de Profesorado y Licenciatura en Educación Inicial y Parvularia, ganadora de movilidad académica en Cuba" href="http://www.uees.edu.sv/?news=estudiante-profesorado-licenciatura-educacion-inicial-parvularia-ganadora-movilidad-academica-cuba "><img width="1024" height="620" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/cuba6.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/02/cuba6.jpg 1024w, http://www.uees.edu.sv/wp-content/uploads/2018/02/cuba6-300x182.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2018/02/cuba6-768x465.jpg 768w" sizes="(max-width: 1024px) 100vw, 1024px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="Estudiante de Profesorado y Licenciatura en Educación Inicial y Parvularia, ganadora de movilidad académica en Cuba" href="http://www.uees.edu.sv/?news=estudiante-profesorado-licenciatura-educacion-inicial-parvularia-ganadora-movilidad-academica-cuba ">Estudiante de Profesorado y Licenciatura en Educación Inicial y Parvularia, ganadora de movilidad académica en Cuba</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="Estudiante de Profesorado y Licenciatura en Educación Inicial y Parvularia, ganadora de movilidad académica en Cuba" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/cuba6.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=estudiante-profesorado-licenciatura-educacion-inicial-parvularia-ganadora-movilidad-academica-cuba" title="Estudiante de Profesorado y Licenciatura en Educación Inicial y Parvularia, ganadora de movilidad académica en Cuba">Details</a></div></div></div></article><!-- .hentry --><article class="post-20780 news type-news status-publish has-post-thumbnail hentry"><div class="image-area"><a title="AFP CRECER PREMIA A 36 EMPRESAS POR CALIDAD Y PAGO PUNTUAL DE COTIZACIONES" href="http://www.uees.edu.sv/?news=afp-crecer-premia-36-empresas-calidad-pago-puntual-cotizaciones "><img width="735" height="468" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/EDH20180216NEG055P_3.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/02/EDH20180216NEG055P_3.jpg 735w, http://www.uees.edu.sv/wp-content/uploads/2018/02/EDH20180216NEG055P_3-300x191.jpg 300w" sizes="(max-width: 735px) 100vw, 735px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="AFP CRECER PREMIA A 36 EMPRESAS POR CALIDAD Y PAGO PUNTUAL DE COTIZACIONES" href="http://www.uees.edu.sv/?news=afp-crecer-premia-36-empresas-calidad-pago-puntual-cotizaciones ">AFP CRECER PREMIA A 36 EMPRESAS POR CALIDAD Y PAGO PUNTUAL DE COTIZACIONES</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="AFP CRECER PREMIA A 36 EMPRESAS POR CALIDAD Y PAGO PUNTUAL DE COTIZACIONES" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/EDH20180216NEG055P_3.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=afp-crecer-premia-36-empresas-calidad-pago-puntual-cotizaciones" title="AFP CRECER PREMIA A 36 EMPRESAS POR CALIDAD Y PAGO PUNTUAL DE COTIZACIONES">Details</a></div></div></div></article><!-- .hentry --><article class="post-20768 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2018"><div class="image-area"><a title="FACULTAD DE ODONTOLOGÍA ESTUDIANTES DEL TAO, RECIBIERON TALLER DE GLOBOFLEXIA" href="http://www.uees.edu.sv/?news=facultad-odontologia-estudiantes-del-tao-recibieron-taller-globoflexia "><img width="1024" height="507" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/globoportada.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/02/globoportada.jpg 1024w, http://www.uees.edu.sv/wp-content/uploads/2018/02/globoportada-300x149.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2018/02/globoportada-768x380.jpg 768w" sizes="(max-width: 1024px) 100vw, 1024px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="FACULTAD DE ODONTOLOGÍA ESTUDIANTES DEL TAO, RECIBIERON TALLER DE GLOBOFLEXIA" href="http://www.uees.edu.sv/?news=facultad-odontologia-estudiantes-del-tao-recibieron-taller-globoflexia ">FACULTAD DE ODONTOLOGÍA ESTUDIANTES DEL TAO, RECIBIERON TALLER DE GLOBOFLEXIA</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="FACULTAD DE ODONTOLOGÍA ESTUDIANTES DEL TAO, RECIBIERON TALLER DE GLOBOFLEXIA" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/globoportada.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=facultad-odontologia-estudiantes-del-tao-recibieron-taller-globoflexia" title="FACULTAD DE ODONTOLOGÍA ESTUDIANTES DEL TAO, RECIBIERON TALLER DE GLOBOFLEXIA">Details</a></div></div></div></article><!-- .hentry --><article class="post-20659 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2018"><div class="image-area"><a title="VICERRECTORÍA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL REUNIÓN GENERAL PROGRAMA BECAS UEES" href="http://www.uees.edu.sv/?news=vicerrectoria-investigacion-proyeccion-social-reunion-general-programa-becas-uees "><img width="1000" height="573" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/foto5-e1520886737931.jpg" class="thumbnail wp-post-image" alt="" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="VICERRECTORÍA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL REUNIÓN GENERAL PROGRAMA BECAS UEES" href="http://www.uees.edu.sv/?news=vicerrectoria-investigacion-proyeccion-social-reunion-general-programa-becas-uees ">VICERRECTORÍA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL REUNIÓN GENERAL PROGRAMA BECAS UEES</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="VICERRECTORÍA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL REUNIÓN GENERAL PROGRAMA BECAS UEES" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/foto5-e1520886737931.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=vicerrectoria-investigacion-proyeccion-social-reunion-general-programa-becas-uees" title="VICERRECTORÍA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL REUNIÓN GENERAL PROGRAMA BECAS UEES">Details</a></div></div></div></article><!-- .hentry --><article class="post-20655 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2018"><div class="image-area"><a title="INAUGURACIÓN CICLO ACADÉMICO 01-2018 Y FOOD COURT UEES" href="http://www.uees.edu.sv/?news=inauguracion-ciclo-academico-01-2018-food-court-uees "><img width="800" height="434" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/foto1.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/02/foto1.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2018/02/foto1-300x163.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2018/02/foto1-768x417.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="INAUGURACIÓN CICLO ACADÉMICO 01-2018 Y FOOD COURT UEES" href="http://www.uees.edu.sv/?news=inauguracion-ciclo-academico-01-2018-food-court-uees ">INAUGURACIÓN CICLO ACADÉMICO 01-2018 Y FOOD COURT UEES</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="INAUGURACIÓN CICLO ACADÉMICO 01-2018 Y FOOD COURT UEES" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/foto1.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=inauguracion-ciclo-academico-01-2018-food-court-uees" title="INAUGURACIÓN CICLO ACADÉMICO 01-2018 Y FOOD COURT UEES">Details</a></div></div></div></article><!-- .hentry --><article class="post-20533 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2018"><div class="image-area"><a title="FACULTAD DE INGENIERÍAS &#8211; FIRMA DE CARTA DE ENTENDIMIENTO CON LA SECRETARÍA DE PARTICIPACIÓN, TRANSPARENCIA Y ANTICORRUPCIÓN" href="http://www.uees.edu.sv/?news=firma-carta-entendimiento-la-secretaria-participacion-transparencia-anticorrupcion "><img width="900" height="528" src="http://www.uees.edu.sv/wp-content/uploads/2018/02/carta4.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2018/02/carta4.jpg 900w, http://www.uees.edu.sv/wp-content/uploads/2018/02/carta4-300x176.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2018/02/carta4-768x451.jpg 768w" sizes="(max-width: 900px) 100vw, 900px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="FACULTAD DE INGENIERÍAS &#8211; FIRMA DE CARTA DE ENTENDIMIENTO CON LA SECRETARÍA DE PARTICIPACIÓN, TRANSPARENCIA Y ANTICORRUPCIÓN" href="http://www.uees.edu.sv/?news=firma-carta-entendimiento-la-secretaria-participacion-transparencia-anticorrupcion ">FACULTAD DE INGENIERÍAS &#8211; FIRMA DE CARTA DE ENTENDIMIENTO CON LA SECRETARÍA DE PARTICIPACIÓN, TRANSPARENCIA Y ANTICORRUPCIÓN</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="FACULTAD DE INGENIERÍAS &#8211; FIRMA DE CARTA DE ENTENDIMIENTO CON LA SECRETARÍA DE PARTICIPACIÓN, TRANSPARENCIA Y ANTICORRUPCIÓN" href="http://www.uees.edu.sv/wp-content/uploads/2018/02/carta4.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=firma-carta-entendimiento-la-secretaria-participacion-transparencia-anticorrupcion" title="FACULTAD DE INGENIERÍAS &#8211; FIRMA DE CARTA DE ENTENDIMIENTO CON LA SECRETARÍA DE PARTICIPACIÓN, TRANSPARENCIA Y ANTICORRUPCIÓN">Details</a></div></div></div></article><!-- .hentry --></div></div><!-- carousel-container --></div><!-- carousel-wrap --></div></div><div id="panel-14611-1-0-2" class="so-panel widget widget_mo-post-snippets-carousel panel-last-child" data-index="4" ><div class="so-widget-mo-post-snippets-carousel so-widget-mo-post-snippets-carousel-default-d75171398898"><script type="text/javascript">
jQuery(document).ready(function($) {jQuery('#news-carousel .slides').owlCarousel({navigation: false,navigationText: ["<i class=\"icon-uniF489\"></i>","<i class=\"icon-uniF488\"></i>"],scrollPerPage: false,items: 4,itemsDesktop: [1199,4],itemsDesktopSmall: [979,5],itemsTablet: [768,4],itemsTabletSmall: [640,2],itemsMobile: [479,1],autoPlay: 5000,stopOnHover: true,pagination: false,rewindSpeed: 200,slideSpeed: 800,paginationSpeed: "0"})});
</script>
<div class="carousel-wrap"><div id ="news-carousel" class="carousel-container"><div class="slides image-grid post-snippets  owl-carousel"><article class="post-11831 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE INGENIERÍAS CLAUSURA DEL PROGRAMA: “NIÑOS TALENTOS EN TECNOLOGÍAS DE INFORMACIÓN Y LA COMUNICACIÓN 2017”" href="http://www.uees.edu.sv/?news=library-reopens-post-renovation "><img width="800" height="510" src="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia6.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia6.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia6-300x191.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia6-768x490.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE INGENIERÍAS CLAUSURA DEL PROGRAMA: “NIÑOS TALENTOS EN TECNOLOGÍAS DE INFORMACIÓN Y LA COMUNICACIÓN 2017”" href="http://www.uees.edu.sv/?news=library-reopens-post-renovation ">UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE INGENIERÍAS CLAUSURA DEL PROGRAMA: “NIÑOS TALENTOS EN TECNOLOGÍAS DE INFORMACIÓN Y LA COMUNICACIÓN 2017”</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE INGENIERÍAS CLAUSURA DEL PROGRAMA: “NIÑOS TALENTOS EN TECNOLOGÍAS DE INFORMACIÓN Y LA COMUNICACIÓN 2017”" href="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia6.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=library-reopens-post-renovation" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE INGENIERÍAS CLAUSURA DEL PROGRAMA: “NIÑOS TALENTOS EN TECNOLOGÍAS DE INFORMACIÓN Y LA COMUNICACIÓN 2017”">Details</a></div></div></div></article><!-- .hentry --><article class="post-12058 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="PROCURADURÍA GENERAL DE LA REPÚBLICA OTORGÓ CERTIFICADO DE ACREDITACIÓN Y FUNCIONAMIENTO PARA CENTRO INTEGRADO DE MEDIACIÓN Y SOCORRO JURÍDICO" href="http://www.uees.edu.sv/?news=sports-meet "><img width="800" height="510" src="http://www.uees.edu.sv/wp-content/uploads/2014/10/noticia7.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/10/noticia7.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2014/10/noticia7-300x191.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/10/noticia7-768x490.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="PROCURADURÍA GENERAL DE LA REPÚBLICA OTORGÓ CERTIFICADO DE ACREDITACIÓN Y FUNCIONAMIENTO PARA CENTRO INTEGRADO DE MEDIACIÓN Y SOCORRO JURÍDICO" href="http://www.uees.edu.sv/?news=sports-meet ">PROCURADURÍA GENERAL DE LA REPÚBLICA OTORGÓ CERTIFICADO DE ACREDITACIÓN Y FUNCIONAMIENTO PARA CENTRO INTEGRADO DE MEDIACIÓN Y SOCORRO JURÍDICO</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="PROCURADURÍA GENERAL DE LA REPÚBLICA OTORGÓ CERTIFICADO DE ACREDITACIÓN Y FUNCIONAMIENTO PARA CENTRO INTEGRADO DE MEDIACIÓN Y SOCORRO JURÍDICO" href="http://www.uees.edu.sv/wp-content/uploads/2014/10/noticia7.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=sports-meet" title="PROCURADURÍA GENERAL DE LA REPÚBLICA OTORGÓ CERTIFICADO DE ACREDITACIÓN Y FUNCIONAMIENTO PARA CENTRO INTEGRADO DE MEDIACIÓN Y SOCORRO JURÍDICO">Details</a></div></div></div></article><!-- .hentry --><article class="post-11403 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL INAUGURACIÓN DE SEMANA CULTURAL 2017 “POR UNA CULTURA MEDIOAMBIENTAL SUSTENTABLE”" href="http://www.uees.edu.sv/?news=412-receive-degrees-at-commencement "><img width="800" height="510" src="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia4.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia4.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia4-300x191.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia4-768x490.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL INAUGURACIÓN DE SEMANA CULTURAL 2017 “POR UNA CULTURA MEDIOAMBIENTAL SUSTENTABLE”" href="http://www.uees.edu.sv/?news=412-receive-degrees-at-commencement ">UNIVERSIDAD EVANGÉLICA DE EL SALVADOR VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL INAUGURACIÓN DE SEMANA CULTURAL 2017 “POR UNA CULTURA MEDIOAMBIENTAL SUSTENTABLE”</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL INAUGURACIÓN DE SEMANA CULTURAL 2017 “POR UNA CULTURA MEDIOAMBIENTAL SUSTENTABLE”" href="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia4.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=412-receive-degrees-at-commencement" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL INAUGURACIÓN DE SEMANA CULTURAL 2017 “POR UNA CULTURA MEDIOAMBIENTAL SUSTENTABLE”">Details</a></div></div></div></article><!-- .hentry --><article class="post-11401 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL UNIDAD DE ARTE, CULTURA Y DEPORTES UEES PARTICIPA EN INAUGURACIÓN DE LOS XXXVI JUEGOS DEPORTIVOS ADUSAL 2017" href="http://www.uees.edu.sv/?news=art-work-of-invent-seniors-on-display-at-art-gallery "><img width="800" height="510" src="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia3.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia3.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia3-300x191.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia3-768x490.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL UNIDAD DE ARTE, CULTURA Y DEPORTES UEES PARTICIPA EN INAUGURACIÓN DE LOS XXXVI JUEGOS DEPORTIVOS ADUSAL 2017" href="http://www.uees.edu.sv/?news=art-work-of-invent-seniors-on-display-at-art-gallery ">VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL UNIDAD DE ARTE, CULTURA Y DEPORTES UEES PARTICIPA EN INAUGURACIÓN DE LOS XXXVI JUEGOS DEPORTIVOS ADUSAL 2017</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL UNIDAD DE ARTE, CULTURA Y DEPORTES UEES PARTICIPA EN INAUGURACIÓN DE LOS XXXVI JUEGOS DEPORTIVOS ADUSAL 2017" href="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia3.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=art-work-of-invent-seniors-on-display-at-art-gallery" title="VICERRECTORIA DE INVESTIGACIÓN Y PROYECCIÓN SOCIAL UNIDAD DE ARTE, CULTURA Y DEPORTES UEES PARTICIPA EN INAUGURACIÓN DE LOS XXXVI JUEGOS DEPORTIVOS ADUSAL 2017">Details</a></div></div></div></article><!-- .hentry --><article class="post-11399 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR  DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL  FIRMA DE CONVENIO UEES-GLOBAL VISION CHRISTIAN SHOOL-FUNDACIÓN VÉRITAS" href="http://www.uees.edu.sv/?news=invent-college-named-green-college "><img width="2000" height="1333" src="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2.jpg 2000w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2-300x200.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2-768x512.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2-1024x682.jpg 1024w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2-272x182.jpg 272w" sizes="(max-width: 2000px) 100vw, 2000px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR  DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL  FIRMA DE CONVENIO UEES-GLOBAL VISION CHRISTIAN SHOOL-FUNDACIÓN VÉRITAS" href="http://www.uees.edu.sv/?news=invent-college-named-green-college ">UNIVERSIDAD EVANGÉLICA DE EL SALVADOR  DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL  FIRMA DE CONVENIO UEES-GLOBAL VISION CHRISTIAN SHOOL-FUNDACIÓN VÉRITAS</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR  DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL  FIRMA DE CONVENIO UEES-GLOBAL VISION CHRISTIAN SHOOL-FUNDACIÓN VÉRITAS" href="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia2.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=invent-college-named-green-college" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR  DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL  FIRMA DE CONVENIO UEES-GLOBAL VISION CHRISTIAN SHOOL-FUNDACIÓN VÉRITAS">Details</a></div></div></div></article><!-- .hentry --><article class="post-11397 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="OCTOGÉSIMA CUARTA GRADUACIÓN DE PROFESIONALES UEES ABRIL 2017" href="http://www.uees.edu.sv/?news=invent-student-paper-first-in-scholastic-awards "><img width="2000" height="1333" src="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1.jpg 2000w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1-300x200.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1-768x512.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1-1024x682.jpg 1024w, http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1-272x182.jpg 272w" sizes="(max-width: 2000px) 100vw, 2000px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="OCTOGÉSIMA CUARTA GRADUACIÓN DE PROFESIONALES UEES ABRIL 2017" href="http://www.uees.edu.sv/?news=invent-student-paper-first-in-scholastic-awards ">OCTOGÉSIMA CUARTA GRADUACIÓN DE PROFESIONALES UEES ABRIL 2017</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="OCTOGÉSIMA CUARTA GRADUACIÓN DE PROFESIONALES UEES ABRIL 2017" href="http://www.uees.edu.sv/wp-content/uploads/2014/05/noticia1.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=invent-student-paper-first-in-scholastic-awards" title="OCTOGÉSIMA CUARTA GRADUACIÓN DE PROFESIONALES UEES ABRIL 2017">Details</a></div></div></div></article><!-- .hentry --><article class="post-11409 news type-news status-publish has-post-thumbnail hentry news_category-noticias-2017"><div class="image-area"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE ODONTOLOGÍA-DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL. “FIRMA DE CONVENIO UEES-FEDEX PABLO TESAK”" href="http://www.uees.edu.sv/?news=invent-college-to-celebrate-commencement-on-may-15 "><img width="800" height="510" src="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia5.jpg" class="thumbnail wp-post-image" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia5.jpg 800w, http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia5-300x191.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia5-768x490.jpg 768w" sizes="(max-width: 800px) 100vw, 800px" /></a><div class="image-overlay"></div><div class="image-info"><h4 class="post-title"><a title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE ODONTOLOGÍA-DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL. “FIRMA DE CONVENIO UEES-FEDEX PABLO TESAK”" href="http://www.uees.edu.sv/?news=invent-college-to-celebrate-commencement-on-may-15 ">UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE ODONTOLOGÍA-DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL. “FIRMA DE CONVENIO UEES-FEDEX PABLO TESAK”</a></h4><div class="image-info-buttons"><a class="lightbox-link button transparent" data-gal="prettyPhoto[]" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE ODONTOLOGÍA-DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL. “FIRMA DE CONVENIO UEES-FEDEX PABLO TESAK”" href="http://www.uees.edu.sv/wp-content/uploads/2014/06/noticia5.jpg ">Expand</a><a class="post-link button transparent" href="http://www.uees.edu.sv/?news=invent-college-to-celebrate-commencement-on-may-15" title="UNIVERSIDAD EVANGÉLICA DE EL SALVADOR FACULTAD DE ODONTOLOGÍA-DIRECCIÓN DE RELACIONES Y COOPERACIÓN INTERNACIONAL. “FIRMA DE CONVENIO UEES-FEDEX PABLO TESAK”">Details</a></div></div></div></article><!-- .hentry --></div></div><!-- carousel-container --></div><!-- carousel-wrap --></div></div></div></div></div><div id="pg-14611-2"  class="panel-grid panel-has-style" ><div class="siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-2" data-stretch-type="full-stretched" ><div id="pgc-14611-2-0"  class="panel-grid-cell" ><div id="panel-14611-2-0-0" class="so-panel widget widget_mo-heading panel-first-child" data-index="5" ><div class="so-widget-mo-heading so-widget-mo-heading-default-d75171398898">
<div class="heading1 separator"><h3 class="title"><br /><br />VIDEO INSTITUCIONAL</h3></div></div></div><div id="panel-14611-2-0-1" class="so-panel widget widget_sow-editor panel-last-child" data-index="6" ><div class="so-widget-sow-editor so-widget-sow-editor-base">
<div class="siteorigin-widget-tinymce textwidget">
	<p><iframe width="560" height="315" src="https://www.youtube.com/embed/QKvL8ZyI9EM?rel=0&amp;controls=0&amp;showinfo=0&amp;start=3" frameborder="0" allow="autoplay; encrypted-media" allowfullscreen></iframe></p>
</div>
</div></div></div></div></div><div id="pg-14611-3"  class="panel-grid panel-has-style" ><div class="siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-3" data-stretch-type="full-stretched" ><div id="pgc-14611-3-0"  class="panel-grid-cell" ><div id="panel-14611-3-0-0" class="so-panel widget widget_mo-heading panel-first-child" data-index="7" ><div class="so-widget-mo-heading so-widget-mo-heading-default-d75171398898">
<div class="heading1 separator"><h3 class="title"><br /><br />UNIVERSIDAD EN MOVIMIENTO</h3></div></div></div><div id="panel-14611-3-0-1" class="so-panel widget widget_sow-editor panel-last-child" data-index="8" ><div class="so-widget-sow-editor so-widget-sow-editor-base">
<div class="siteorigin-widget-tinymce textwidget">
	<div class="vc_row wpb_row vc_row-fluid">
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_bounceInDown bounceInDown">
<h2 class="wpb_heading wpb_singleimage_heading">RELACIONES INTERNACIONALES</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=18304" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="194" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/internacional-300x194.jpg" class="vc_single_image-img attachment-medium" alt="" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_bounceInLeft bounceInLeft">
<h2 class="wpb_heading wpb_singleimage_heading">DIRECCIÓN DE INVESTIGACIÓN</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=16411" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="188" src="http://www.uees.edu.sv/wp-content/uploads/2014/10/investigacion3-300x188.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2014/10/investigacion3-300x188.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2014/10/investigacion3-768x480.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2014/10/investigacion3-1024x640.jpg 1024w, http://www.uees.edu.sv/wp-content/uploads/2014/10/investigacion3.jpg 1200w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_bounceInRight bounceInRight">
<h2 class="wpb_heading wpb_singleimage_heading">DIRECCIÓN DE PUBLICACIONES</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=17683" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="194" src="http://www.uees.edu.sv/wp-content/uploads/2017/10/libros111-300x194-1-300x194.jpg" class="vc_single_image-img attachment-medium" alt="" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_bounceInUp bounceInUp">
<h2 class="wpb_heading wpb_singleimage_heading">PROYECCIÓN<br />
 SOCIAL</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=326" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="194" src="http://www.uees.edu.sv/wp-content/uploads/2017/10/proyectosocial_cultura55-300x194.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2017/10/proyectosocial_cultura55-300x194.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2017/10/proyectosocial_cultura55.jpg 700w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
</div>
<div class="vc_row wpb_row vc_row-fluid">
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_rotateIn rotateIn">
<h2 class="wpb_heading wpb_singleimage_heading">CAMPUS UEES</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=135" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="199" src="http://www.uees.edu.sv/wp-content/uploads/2017/04/foto10-300x199.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2017/04/foto10-300x199.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2017/04/foto10-768x510.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2017/04/foto10.jpg 1024w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_fadeInDownBig fadeInDownBig">
<h2 class="wpb_heading wpb_singleimage_heading">ARTE Y CULTURA</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=18294" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="189" src="http://www.uees.edu.sv/wp-content/uploads/2017/04/arte-300x189.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2017/04/arte-300x189.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2017/04/arte-768x483.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2017/04/arte.jpg 960w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_fadeInRightBig fadeInRightBig">
<h2 class="wpb_heading wpb_singleimage_heading">GRADUADOS</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=16448" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="183" src="http://www.uees.edu.sv/wp-content/uploads/2017/04/graduados-300x183.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2017/04/graduados-300x183.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2017/04/graduados-768x467.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2017/04/graduados.jpg 1024w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
<div class="wpb_column vc_column_container vc_col-sm-3">
<div class="vc_column-inner ">
<div class="wpb_wrapper">
<div  class="wpb_single_image wpb_content_element vc_align_center  wpb_animate_when_almost_visible wpb_slideInRight slideInRight">
<h2 class="wpb_heading wpb_singleimage_heading">DEPORTES</h2>
<figure class="wpb_wrapper vc_figure">
			<a href="http://www.uees.edu.sv/?page_id=18290" target="_self" class="vc_single_image-wrapper vc_box_shadow_3d  vc_box_border_grey"><img width="300" height="189" src="http://www.uees.edu.sv/wp-content/uploads/2017/04/baske2m-300x189.jpg" class="vc_single_image-img attachment-medium" alt="" srcset="http://www.uees.edu.sv/wp-content/uploads/2017/04/baske2m-300x189.jpg 300w, http://www.uees.edu.sv/wp-content/uploads/2017/04/baske2m-768x484.jpg 768w, http://www.uees.edu.sv/wp-content/uploads/2017/04/baske2m.jpg 1007w" sizes="(max-width: 300px) 100vw, 300px" /></a><br />
		</figure>
</p></div>
</div>
</div>
</div>
</div>
</div>
</div></div></div></div></div><div id="pg-14611-4"  class="panel-grid panel-has-style" ><div class="siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-4" data-stretch-type="full" id="stats-section" ><div id="pgc-14611-4-0"  class="panel-grid-cell panel-grid-cell-empty" ></div></div></div><div id="pg-14611-5"  class="panel-grid panel-has-style" ><div class="siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-5" data-stretch-type="full-stretched" ><div id="pgc-14611-5-0"  class="panel-grid-cell" ><div id="panel-14611-5-0-0" class="so-panel widget widget_mo-hero-section panel-first-child panel-last-child" data-index="9" ><div class="so-widget-mo-hero-section so-widget-mo-hero-section-default-d75171398898"><div  data-parallax-speed="0.4" class="segment clearfix quote-banner parallax-background parallax-banner"  style="background-image:url(http://www.uees.edu.sv/wp-content/uploads/2016/03/visionymision2.jpg); background-color:#2a9dd6;background-attachment:fixed;"><div class="segment-content"><h2>MISIÓN</h2><div class="text"><p>“Formar profesionales con excelencia académica, conscientes del servicio a sus semejantes y con una ética cristiana basada en las sagradas escrituras para responder a las necesidades y cambios de la sociedad”.</p></div><h2>VISIÓN</h2><div class="text"><p>“Ser la institución de educación superior, líder regional por su excelencia académica e innovación científica y tecnológica; reconocida por su naturaleza y práctica cristiana.”</p></div></div></div><!-- .segment--></div></div></div></div></div><div id="pg-14611-6"  class="panel-grid panel-has-style" ><div class="siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-6" data-stretch-type="full" id="featured-sources" ><div id="pgc-14611-6-0"  class="panel-grid-cell" ><div id="panel-14611-6-0-0" class="so-panel widget widget_mo-heading panel-first-child" data-index="10" ><div class="so-widget-mo-heading so-widget-mo-heading-default-d75171398898">
<div class="heading1 separator"><h3 class="title"><br /><br /><strong>AFILIACIONES</strong></h3></div></div></div><div id="panel-14611-6-0-1" class="so-panel widget widget_sow-editor panel-last-child" data-index="11" ><div class="so-widget-sow-editor so-widget-sow-editor-base">
<div class="siteorigin-widget-tinymce textwidget">
	<p><strong> </strong></p>
<p><strong> </strong></p>
<table style="height: 178px;" border="0" width="750" cellspacing="10" cellpadding="0" align="center">
<tbody>
<tr>
<td align="center" width="127"><img class=" wp-image-16622 aligncenter" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio3.png" alt="" width="127" height="127" /></td>
<td align="center" width="127"><strong><img class="alignnone wp-image-18872 " src="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio44-1.png" alt="" width="126" height="126" /></strong></td>
<td align="center" width="121"><img class=" wp-image-16620 aligncenter" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio1.png" alt="" width="121" height="121" /></td>
<td align="center" width="126"><strong><img class=" wp-image-16621 aligncenter" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/logoconvenio2.png" alt="" width="125" height="125" /></strong></td>
<td align="center" width="189"><img class="alignnone size-full wp-image-19491" src="http://www.uees.edu.sv/wp-content/uploads/2016/03/logopanalExok.png" alt="" width="178" height="151" /></td>
</tr>
</tbody>
</table>
</div>
</div></div></div></div></div><div id="pg-14611-7"  class="panel-grid panel-has-style" ><div class="call-to-action clearfix siteorigin-panels-stretch panel-row-style panel-row-style-for-14611-7" data-stretch-type="full-stretched" ><div id="pgc-14611-7-0"  class="panel-grid-cell panel-grid-cell-empty" ></div></div></div></div>
                        
                    </div>
                    <!-- .entry-content -->

                    
                </article><!-- .hentry -->

                
                
                
                
            
        
        
    </div><!-- #content -->


    </div> <!-- #one-column-template -->


</div><!-- #main .inner -->


</div><!-- #main -->

    
    <footer id="footer">

        <div class="inner">

            
            <div id="sidebars-footer" class="clearfix">

                <div id="sidebar-footer1" class="sidebar clearfix fourcol"><aside id="nav_menu-9" class="widget widget_nav_menu widget-widget_nav_menu"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>Sitios de Interes</span></h3><div class="menu-sitios-de-interes-container"><ul id="menu-sitios-de-interes" class="menu"><li id="menu-item-17751" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17751"><a href="http://www.uees.edu.sv/?page_id=15989">Portal del Estudiante</a></li>
<li id="menu-item-17750" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17750"><a href="http://www.uees.edu.sv/?page_id=322">Portal del Docente</a></li>
<li id="menu-item-17759" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17759"><a href="http://www.uees.edu.sv/?page_id=16503">Biblioteca</a></li>
<li id="menu-item-17744" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17744"><a href="http://www.uees.edu.sv/?page_id=17683">Editorial UEES</a></li>
<li id="menu-item-17746" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17746"><a href="http://www.uees.edu.sv/?page_id=16151">Escuela de Posgrado</a></li>
<li id="menu-item-17745" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17745"><a href="http://www.uees.edu.sv/?page_id=16237">EPOUEES</a></li>
<li id="menu-item-17755" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17755"><a href="http://www.uees.edu.sv/?page_id=17694">Cursos</a></li>
<li id="menu-item-17757" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17757"><a href="http://www.uees.edu.sv/?page_id=16448">Graduados</a></li>
<li id="menu-item-17758" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17758"><a href="http://www.uees.edu.sv/?page_id=14242">UEES Virtual</a></li>
</ul></div></div></aside><aside id="nav_menu-8" class="widget widget_nav_menu widget-widget_nav_menu"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>Facultades</span></h3><div class="menu-facultades-container"><ul id="menu-facultades" class="menu"><li id="menu-item-17764" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17764"><a href="http://www.uees.edu.sv/?page_id=15566">Facultad de Medicina</a></li>
<li id="menu-item-17765" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17765"><a href="http://www.uees.edu.sv/?page_id=15588">Facultad de Odontología</a></li>
<li id="menu-item-17760" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17760"><a href="http://www.uees.edu.sv/?page_id=15709">Facultad de Ciencias Jurídicas</a></li>
<li id="menu-item-17761" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17761"><a href="http://www.uees.edu.sv/?page_id=15758">Facultad de Ciencias Sociales</a></li>
<li id="menu-item-17762" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17762"><a href="http://www.uees.edu.sv/?page_id=15892">Facultad de Ciencias Empresariales y Económicas</a></li>
<li id="menu-item-17763" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-17763"><a href="http://www.uees.edu.sv/?page_id=15691">Facultad de Ingenierías</a></li>
</ul></div></div></aside></div><div id="sidebar-footer2" class="sidebar clearfix fourcol"><aside id="text-12" class="widget widget_text widget-widget_text"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>Contactenos</span></h3>			<div class="textwidget"><div class="frm_forms  with_frm_style frm_style_formidable-style" id="frm_form_3_container" >
<form enctype="multipart/form-data" method="post" class="frm-show-form " id="form_s7lsu"  >
<div class="frm_form_fields ">
<fieldset>
<legend class="frm_screen_reader">Contactenos</legend>

<div class="frm_fields_container">
<input type="hidden" name="frm_action" value="create" />
<input type="hidden" name="form_id" value="3" />
<input type="hidden" name="frm_hide_fields_3" id="frm_hide_fields_3" value="" />
<input type="hidden" name="form_key" value="s7lsu" />
<input type="hidden" name="item_meta[0]" value="" />
<input type="hidden" id="frm_submit_entry_3" name="frm_submit_entry_3" value="89dc5da6c1" /><input type="hidden" name="_wp_http_referer" value="/" /><label for="frm_verify_3" class="frm_screen_reader frm_hidden">If you are human, leave this field blank.</label>
<input type="text" class="frm_hidden frm_verify" id="frm_verify_3" name="frm_verify" value=""  />
<div id="frm_field_11_container" class="frm_form_field form-field  frm_required_field frm_top_container">
    <label for="field_6jl31" class="frm_primary_label">Nombre:
        <span class="frm_required">*</span>
    </label>
    <textarea name="item_meta[11]" id="field_6jl31" rows="1"  style="width:250px" cols="27" data-reqmsg="Este campo no puede estar en blanco." data-invmsg="Nombre: no es válido" class="auto_width"  ></textarea>
    
    
</div>
<div id="frm_field_13_container" class="frm_form_field form-field  frm_required_field frm_top_container">
    <label for="field_n52bl" class="frm_primary_label">Correo electronico
        <span class="frm_required">*</span>
    </label>
    <input type="email" id="field_n52bl" name="item_meta[13]" value=""  style="width:250px" maxlength="50" data-reqmsg="Este campo no puede estar en blanco." data-invmsg="Correo electronico no es válido" class="auto_width"  />
    
    
</div>
<div id="frm_field_14_container" class="frm_form_field form-field  frm_top_container">
    <label for="field_mfh50" class="frm_primary_label">Comentario o Mensaje
        <span class="frm_required"></span>
    </label>
    <textarea name="item_meta[14]" id="field_mfh50" rows="5"  style="width:300px" cols="33" data-invmsg="Comentario o Mensaje no es válido" class="auto_width"  ></textarea>
    
    
</div>
<div id="frm_field_28_container" class="frm_form_field form-field  frm_none_container">
    <label  class="frm_primary_label">reCAPTCHA
        <span class="frm_required"></span>
    </label>
    
    
    
</div>
<input type="hidden" name="item_key" value="" />
<div class="frm_submit">

<button class="frm_button_submit" type="submit"  >Enviar</button>

</div></div>
</fieldset>
</div>
</form>
</div>
</div>
		</div></aside><aside id="text-11" class="widget widget_text widget-widget_text"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>Contador de Visitas</span></h3>			<div class="textwidget"><script type="text/javascript" src="https://counter2.freecounter.ovh/private/counter.js?c=bqkw1hmbxd1qgj2h6sn4clq4xylmz5n3&down=async" async></script>

<noscript></noscript><a title="contador de visitas para tumblr" href="https://www.contadorvisitasgratis.com"><img title="contador de visitas para tumblr" src="https://counter2.freecounter.ovh/private/contadorvisitasgratis.php?c=bqkw1hmbxd1qgj2h6sn4clq4xylmz5n3" alt="contador de visitas para tumblr" border="0" /></a></div>
		</div></aside></div><div id="sidebar-footer3" class="sidebar clearfix fourcol last"><aside id="text-10" class="widget widget_text widget-widget_text"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>UEES</span></h3>			<div class="textwidget"><p>Universidad Evangélica de El Salvador<br />
Prolongación Alameda Juan Pablo II,<br />
Calle  El Carmen, San Antonio Abad,<br />
San Salvador, El Salvador<br />
Conmutador: 2275-4000,<br />
Fax: 2275-4040</p>
</div>
		</div></aside><aside id="sow-image-2" class="widget widget_sow-image widget-widget_sow-image"><div class="widget-wrap widget-inside"><div class="so-widget-sow-image so-widget-sow-image-default-642c5433d908">

<div class="sow-image-container">
	<img src="http://www.uees.edu.sv/wp-content/uploads/2018/01/acreditacion2.jpg" title="Inicio" 		class="so-widget-image"/>
</div>

</div></div></aside><aside id="mo-social-networks-widget-2" class="widget social-networks-widget widget-social-networks-widget"><div class="widget-wrap widget-inside"><h3 class="widget-title"><span>Búscanos en las redes</span></h3><ul class="social-list clearfix"><li><a class="facebook" href="https://www.facebook.com/ueesoficial/" target="_blank" title="Follow on Facebook"><i class="icon-facebook8"></i></a></li><li><a class="twitter" href="https://twitter.com/ueesoficial" target="_blank" title="Subscribe to Twitter Feed"><i class="icon-twitter2"></i></a></li><li><a class="youtube" href="https://www.youtube.com/channel/UCZ3m1ZKVzbsyuB3ZZlgXegA" target="_blank" title="Subscribe to the YouTube channel"><i class="icon-youtube4"></i></a></li><li><a class="instagram" href="https://www.instagram.com/explore/locations/1012393993/" target="_blank" title="View Instagram Feed"><i class="icon-instagram5"></i></a></li></ul></div></aside><aside id="mo-button-2" class="widget widget_mo-button widget-widget_mo-button"><div class="widget-wrap widget-inside"><div class="so-widget-mo-button so-widget-mo-button-default-d75171398898"><div style="text-align:center;float:center;"><a class= "button  blue rounded" href="https://mail.uees.edu.sv/owa/auth/logon.aspx?replaceCurrent=1&#038;reason=2&#038;url=https%3a%2f%2fmail.uees.edu.sv%2fowa" target="_blank">Correo Institucional</a></div></div></div></aside><aside id="mo-button-3" class="widget widget_mo-button widget-widget_mo-button"><div class="widget-wrap widget-inside"><div class="so-widget-mo-button so-widget-mo-button-default-d75171398898"><div style="text-align:center;float:center;"><a class= "button  blue rounded" href="http://www.uees.edu.sv/pdf/Acceso_OWA.pdf" target="_blank">Manual de Usuario</a></div></div></div></aside></div>
            </div>
            <!-- #sidebars-footer -->

            
        </div>

    </footer> <!-- #footer -->

    

<footer id="footer-bottom">

    <div class="inner">

        
        <div id="footer-bottom-text">Copyright &#169; 2018 <a class="site-link" href="http://www.uees.edu.sv" title="Universidad Evangélica de El Salvador" rel="home"><span>Universidad Evangélica de El Salvador</span></a>. Powered by <a class="wp-link" href="http://wordpress.org" title="Powered by WordPress"><span>WordPress</span></a> and <a class="theme-link" href="" title="Invent"><span>Invent</span></a></div>
        <a id="go-to-top" href="#" title="Back to top">Go Top</a>
    </div>

</footer><!-- #footer-bottom -->

</div><!-- #container -->


<div class="hidden"><script type="text/javascript">

  var _gaq = _gaq || [];
  _gaq.push(['_setAccount', 'UA-33010281-1']);
  _gaq.push(['_trackPageview']);

  (function() {
    var ga = document.createElement('script'); ga.type = 'text/javascript'; ga.async = true;
    ga.src = ('https:' == document.location.protocol ? 'https://ssl' : 'http://www') + '.google-analytics.com/ga.js';
    var s = document.getElementsByTagName('script')[0]; s.parentNode.insertBefore(ga, s);
  })();

</script></div>		<script type="text/javascript">
			function revslider_showDoubleJqueryError(sliderID) {
				var errorMessage = "Revolution Slider Error: You have some jquery.js library include that comes after the revolution files js include.";
				errorMessage += "<br> This includes make eliminates the revolution slider libraries, and make it not work.";
				errorMessage += "<br><br> To fix it you can:<br>&nbsp;&nbsp;&nbsp; 1. In the Slider Settings -> Troubleshooting set option:  <strong><b>Put JS Includes To Body</b></strong> option to true.";
				errorMessage += "<br>&nbsp;&nbsp;&nbsp; 2. Find the double jquery.js include and remove it.";
				errorMessage = "<span style='font-size:16px;color:#BC0C06;'>" + errorMessage + "</span>";
					jQuery(sliderID).show().html(errorMessage);
			}
		</script>
		<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/livemesh-siteorigin-widgets/assets/js/modernizr-custom.min.js?ver=1.7.3'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/livemesh-siteorigin-widgets/assets/js/jquery.waypoints.min.js?ver=1.7.3'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var lsow_settings = {"mobile_width":"780","custom_css":""};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/livemesh-siteorigin-widgets/assets/js/lsow-frontend.min.js?ver=1.7.3'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.tools.min.js?ver=1.2.7'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.validate.min.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/drop-downs.js?ver=1.4.8'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/waypoints.js?ver=2.0.2'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.plugins.lib.js?ver=1.0'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/skrollr.min.js?ver=1.0'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.mb.YTPlayer.js?ver=1.0'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.flexslider.js?ver=1.2'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/owl.carousel.min.js?ver=4.1'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/jquery.prettyPhoto.js?ver=3.1.6'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/isotope/dist/isotope.pkgd.min.js?ver=5.2'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/imagesloaded.pkgd.min.js?ver=4.1.1'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-includes/js/comment-reply.min.js?ver=4.7.5'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/slider.js?ver=1.0'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var mo_theme = {"name_required":"Please provide your name","name_format":"Your name must consist of at least 5 characters","email_required":"Please provide a valid email address","url_required":"Please provide a valid URL","phone_required":"Minimum 5 characters required","message_required":"Please input the message","message_format":"Your message must be at least 15 characters long","success_message":"Your message has been sent. Thanks!","blog_url":"http:\/\/www.uees.edu.sv","loading_portfolio":"Loading the next set of posts...","finished_loading":"No more items to load..."};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/main.js?ver=1.0'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-includes/js/hoverIntent.min.js?ver=1.8.1'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var megamenu = {"timeout":"300","interval":"100"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/megamenu/js/maxmegamenu.js?ver=2.4.1.5'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/js/dist/js_composer_front.min.js?ver=5.2'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/js_composer/assets/lib/waypoints/waypoints.min.js?ver=5.2'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-includes/js/wp-embed.min.js?ver=4.7.5'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var frm_js = {"ajax_url":"http:\/\/www.uees.edu.sv\/wp-admin\/admin-ajax.php","images_url":"http:\/\/www.uees.edu.sv\/wp-content\/plugins\/formidable\/images","loading":"Loading\u2026","remove":"Eliminar","offset":"4","nonce":"9e032c9dbb","id":"ID","no_results":"Ninguna resultado coincide","file_spam":"That file looks like Spam.","empty_fields":"Please complete the preceding required fields before uploading a file."};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/plugins/formidable/js/frm.min.js?ver=3.0.06'></script>
<script type='text/javascript' defer="defer" async="async" src='https://www.google.com/recaptcha/api.js?onload=frmRecaptcha&#038;render=explicit&#038;hl=es&#038;ver=4.7.5'></script>
<script type='text/javascript' src='http://www.uees.edu.sv/wp-content/themes/invent5/js/libs/waypoints.sticky.min.js?ver=2.0.2'></script>
<script type="text/javascript">document.body.className = document.body.className.replace("siteorigin-panels-before-js","");</script>
</body>
</html>