
<html xmlns="http://www.w3.org/1999/xhtml"
      xmlns:og="http://ogp.me/ns#"
      xmlns:fb="https://www.facebook.com/2008/fbml">  

    <head>
	    
	    <!-- Start Alexa Certify Javascript -->
<script type="text/javascript">
_atrk_opts = { atrk_acct:"jCMMm1a4KM+2cv", domain:"lapagina.com.sv",dynamic: true};
(function() { var as = document.createElement('script'); as.type = 'text/javascript'; as.async = true; as.src = "https://d31qbv1cthcecs.cloudfront.net/atrk.js"; var s = document.getElementsByTagName('script')[0];s.parentNode.insertBefore(as, s); })();
</script>
<noscript><img src="https://d5nxst8fruw4z.cloudfront.net/atrk.gif?account=jCMMm1a4KM+2cv" style="display:none" height="1" width="1" alt="" /></noscript>
<!-- End Alexa Certify Javascript -->  

<script>
  (function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
  (i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
  m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
  })(window,document,'script','//www.google-analytics.com/analytics.js','ga');

  ga('create', 'UA-72603819-1', 'auto');
  ga('send', 'pageview');
  

</script>
		<link rel="icon" href="http://www.lapagina.com.sv/favicon.ico" type="image/x-icon" />
		<link rel="shortcut icon" href="http://lapagina.com.sv/favicon.ico" type="image/x-icon" />
        <meta http-equiv="Content-Type" content="text/html; charset=ISO-8859-1" />




        
        <title>Diario digital de noticias de El Salvador</title>
        <meta name="title" content="Diario digital de noticias de El Salvador" />
        <meta name="DC.Title" content="Diario digital de noticias de El Salvador" />
        <meta http-equiv="title" content="Diario digital de noticias de El Salvador" />
        <meta name="Keywords" content="Diario digital de actualidad de El Salvador, noticias El Salvador, informaciÛn El Salvador, polÌtica El Salvador, deportes El Salvador, Jet set El Salvador" />
        <meta http-equiv="keywords" content="Diario digital de actualidad de El Salvador, noticias El Salvador, informaciÛn El Salvador, polÌtica El Salvador, deportes El Salvador, Jet set El Salvador" />
        	                <meta name="Description" content="Noticias y actualidad de El Salvador. Informaci�n y opini�n sobre pol�tica, deportes y sociedad en el Salvador" />
            <meta http-equiv="description" content="Noticias y actualidad de El Salvador. Informaci�n y opini�n sobre pol�tica, deportes y sociedad en el Salvador" />
            <meta http-equiv="DC.Description" content="Noticias y actualidad de El Salvador. Informaci�n y opini�n sobre pol�tica, deportes y sociedad en el Salvador" />
                <meta name="author" content="Peri�dico Digital La P�gina" />
        <meta name="DC.Creator" content="Peri�dico Digital La P�gina" />
        <meta name="vw96.objectype" content="Homepage" />
        <meta name="resource-type" content="Homepage" />
        <meta name="distribution" content="all" />
        <meta name="robots" content="all" />
        <meta name="language" content="es" />
        <meta http-equiv="Refresh" content="900">
   
        <link href="/estilos/general.css?v=1.55" rel="stylesheet" type="text/css" />
        <link href="/estilos/contenidos.css" rel="stylesheet" type="text/css" />
        <link rel="stylesheet" href="https://maxcdn.bootstrapcdn.com/font-awesome/4.5.0/css/font-awesome.min.css">
		<link rel="stylesheet" href="/social/css/social-share-kit.css" type="text/css">
		
        <script type='text/javascript' src='/js/funciones.js'></script>
        
        <script type='text/javascript' src='/js/js_st.js'></script>
        <ins data-revive-zoneid="1492" data-revive-id="1cc6fd924369584af6e3764ee37b0e18"></ins>
		<script async src="//ads.latinongroup.com/delivery/asyncjs.php"></script>
        
        <script type='text/javascript' src='https://partner.googleadservices.com/gampad/google_service.js'></script>
        <script type='text/javascript'>
                GS_googleAddAdSenseService("ca-pub-3300961026697968");
                GS_googleEnableAllServices();
        </script>
        <script type='text/javascript'>
                GA_googleAddSlot("ca-pub-3300961026697968", "cabecera_derecha");
                GA_googleAddSlot("ca-pub-3300961026697968", "cabecera_izquierda");
                GA_googleAddSlot("ca-pub-3300961026697968", "footer");
                GA_googleAddSlot("ca-pub-3300961026697968", "footer_centro");
                GA_googleAddSlot("ca-pub-3300961026697968", "footer_derecha");
                GA_googleAddSlot("ca-pub-3300961026697968", "footer_Izq");
                GA_googleAddSlot("ca-pub-3300961026697968", "lateral_derecho_1");
                GA_googleAddSlot("ca-pub-3300961026697968", "lateral_derecho_2");
                GA_googleAddSlot("ca-pub-3300961026697968", "lateral_derecho_3");
                GA_googleAddSlot("ca-pub-3300961026697968", "lateral_derecho_4");
                GA_googleAddSlot("ca-pub-3300961026697968", "lateral_derecho_5");
                GA_googleAddSlot("ca-pub-3300961026697968", "Notas_bottom");                
        </script>
        
        <script type='text/javascript'>
                GA_googleFetchAds();
        </script>
        

    </head>
<script type="text/javascript" src="//s7.addthis.com/js/300/addthis_widget.js#pubid=ra-56c2c3254bcb587c" async="async"></script>


    <body>
		<div id="base_header">
            <div id="banners_top">
                <table width="967" border="0" cellpadding="0" cellspacing="0">
                    <tr>
                        <td>
                            <div class="contenedor_banner">
                                <!-- cabecera_izquierda -->
                                <script type='text/javascript'>
                                        GA_googleFillSlot("cabecera_izquierda");
                                </script>
                            </div>
                        </td>
                        <td>
                            <!-- cabecera_derecha -->
                            <div class="contenedor_banner">
                                <script type='text/javascript'>
                                        GA_googleFillSlot("cabecera_derecha");
                                </script>
                            </div>
                        </td>
                    </tr>
                </table>
            </div>
            <div id="header">
                <script>
                        function enviar_busqueda_cab(){
                            document.getElementById("form_cab").submit();
                        }
                </script>
                <form id="form_cab" action="http://www.lapagina.com.sv/res_busqueda.php" method="POST"><input type="hidden" name="pag" value="1">
                        <table width="995" border="0" cellpadding="0" cellspacing="0">
                            <tr>
                                <td><table width="995" border="0" cellpadding="0" cellspacing="0">
                                        <tr>
                                            <td>
                                                <a href="http://www.lapagina.com.sv/">
                                                    <img src="http://www.lapagina.com.sv/images/header/logo_new_.png" border="0" width="501" height="101" />
                                                </a>
                                            </td>
                                            <td valign="bottom"><table width="100%" border="0" cellpadding="0" cellspacing="0">
                                                    <tr>
	                                                    
                                                                                                                <td height="30" class="fecha">

                                                            <div class="ssk_con">
	                                                                 
                                                                <span class="ssk_txt">S&Iacute;GUENOS EN</span>
                                                                <a href="http://fb.me/DiarioLaPaginaSV" target="_blank" class="ssk ssk-facebook" ></a>
																<a href="http://www.twitter.com/lapagina" target="_blank" class="ssk ssk-twitter"></a>
															</div>

                                                            <span style="float: right; margin-top: 25px;">Mi&eacute;rcoles 21 de Marzo de 2018</span>

                                                        </td>
                                                    </tr>
                                                    <tr>
                                                        <td height="40"><table width="100%" border="0" cellpadding="0" cellspacing="0">
                                                                <tr>
                                                                    <td class="linkshd">
	                                                                    <a class="bhead" href="http://www.lapagina.com.sv/boletines.php"><i class="fa fa-paper-plane"></i> boletines</a>
	                                                                    <a class="bhead" href="http://www.lapagina.com.sv/rss.php"><i class="fa fa-rss"></i> RSS</a>
	                                                                    <a class="bhead" href="http://www.lapagina.com.sv/hemeroteca.php"><i class="fa fa-archive"></i> Hemeroteca</a>
	                                                                </td>
                                                                    <td class="searchd" width="210">
	                                                                    <form id="newsearch" method="get" action="javascript:enviar_busqueda_cab()">
		                                                                    <i class="fa fa-search"></i><input type="text" name="buscador" id="buscador" /><input type="submit" value="buscar" class="tfbutton">
	                                                                </td>
                                                                </tr>
                                                            </table></td>
                                                    </tr>
                                                </table></td>
                                        </tr>
                                    </table></td>
                            </tr>
                        </table>
                </form>
            </div>
        </div>
<div class="base_menu">
  <div id="menu_top">
    <p class="botones"><a href="http://www.lapagina.com.sv/portada"  style='color:#ffffff'>PORTADA</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/nacionales" >NACIONALES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/internacionales" >INTERNACIONALES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/entrevistas" >entrevistas</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/empresarial" >empresarial</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/opinion" >OPINI&Oacute;N</a> </p>
    <p class="botones"><a href="http://www.lapagina.com.sv/cultura" >CULTURA</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/deportes" >DEPORTES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/jetset" >JET SET</a></p>
   <p class="boton_fin"><a href="http://www.lapagina.com.sv/curiosidades"  ?>Curiosidades</a></p>
    
  </div>
</div>
		<!---
		<div class="top_especial">
			<a href="http://www.lapagina.com.sv/especiales/resumen2016" target="_self"><img src="images/especiales/resumen_DLP_2016.jpg" border="0"></a>
			
		</div> --->
		
		<div id="base_contenidos" data-sticky_parent>
		  <div id="col_principal">
		    <div id="nota_feat">
		      			   <h3 class="titulo-link"><a href="http://www.lapagina.com.sv/nacionales/137553/2018/03/21/Avianca-suspende-11-vuelos-a-El-Salvador-y-Bogota-por-tormenta-Toby" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Avianca suspende 11 vuelos a El Salvador y Bogot� por tormenta Toby</a></h3>
		      <div class="img_destacada">				
	              <a href="http://www.lapagina.com.sv/nacionales/137553/2018/03/21/Avianca-suspende-11-vuelos-a-El-Salvador-y-Bogota-por-tormenta-Toby"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/JSUA_YXZpb25lcy5qcGc=.jpg" width="" style="margin-bottom:0px;margin-right:5px;" alt=""/></a></div>
		      <div id="texto_notaDestacada">
		        <h1 class="seccion-link"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>   </h1>
		       
		        <div class="desta_cuerpo">
                <p class="desta_lead">La suspensi�n de los vuelos se debe a la tormenta de nieve &ldquo;Toby&rdquo; que azota desde ayer la costa este de los Estados Unidos.
�

</p></div>
		        <div class="div_puntos_pp"></div>
		        		        <div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137553/2018/03/21/Avianca-suspende-11-vuelos-a-El-Salvador-y-Bogota-por-tormenta-Toby#comentarios"> (0) Comentarios</a></div>
		        </div>
		      
		    </div>
		   
		    <div class="div_puntos"></div>
		    <div id="col_01">
		    
		        <div class="name_">LA FRASE</div>
    <div class="frase">
	    <a href="">
        	<div class="img_frase"></div>
			<div class="quote"><p>Esta democracia nueva, joven, necesita que los ciudadanos asuman su compromiso de elegir con el voto secreto		
	</p></div>
			<p class="autor">Salvador S�nchez Cer�n, Presidente de la Rep�blica</p>
	    </a>
    </div>
	  
		      		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137552/2018/03/21/Senalan-conflicto-de-competencias-entre-Sala-de-lo-Civil-y-Juzgado-Especializado-por-caso-diputado-Cardoza"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/QCJQ_ZmlzY2FsX2V4dGluY2lvbl9kZV9kb21pbmlvLmpw.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt="Fiscal Anticorrupci�n, H�ctor Rodr�guez, present� el documento ante la Sala de lo Civil/ Fotograf�a: FGR"/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137552/2018/03/21/Senalan-conflicto-de-competencias-entre-Sala-de-lo-Civil-y-Juzgado-Especializado-por-caso-diputado-Cardoza" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Se�alan conflicto de competencias entre Sala de lo Civil y Juzgado Especializado por caso diputado Cardoza</a></h2>
		      	<p class="texto_nota"> El fiscal Anticorrupci�n pidi� que sea el pleno de la CSJ (los 15 magistrados) quienes resuelvan en el proceso sobre el caso de Reynaldo Cardoza.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137552/2018/03/21/Senalan-conflicto-de-competencias-entre-Sala-de-lo-Civil-y-Juzgado-Especializado-por-caso-diputado-Cardoza#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137546/2018/03/21/Carcel-para-�La-vaca�-y-33-testaferros-de-la-MS-capturados-en-operacion-libertad"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/BRXD_dmFjYS5KUEc=.JPG" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137546/2018/03/21/Carcel-para-�La-vaca�-y-33-testaferros-de-la-MS-capturados-en-operacion-libertad" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">C�rcel para �La vaca� y 33 testaferros de la MS capturados en operaci�n libertad</a></h2>
		      	<p class="texto_nota"> (VIDEO) Los sujetos se encargaban de lavar dinero de la estructura criminal MS que opera en varios municipios del departamento de La Libertad.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137546/2018/03/21/Carcel-para-�La-vaca�-y-33-testaferros-de-la-MS-capturados-en-operacion-libertad#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137544/2018/03/21/Cancilleria-anuncia-datos-preliminares-sobre-el-TPS"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/GKYT_Q2FuY2lsbGVyYXNkYXRwcy5KUEc=.JPG" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137544/2018/03/21/Cancilleria-anuncia-datos-preliminares-sobre-el-TPS" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Canciller�a anuncia datos preliminares sobre el TPS</a></h2>
		      	<p class="texto_nota"> En el marco de la reinscripci�n, el canciller explic� que se retomar�n las gestiones para buscar una alternativa migratoria permanente.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137544/2018/03/21/Cancilleria-anuncia-datos-preliminares-sobre-el-TPS#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137550/2018/03/21/Bomberos-evitan-que-camion-cisterna-explote-con-10-mil-galones-de-combustible"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/UHXO_Ym9tYmVyb3MuanBn.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137550/2018/03/21/Bomberos-evitan-que-camion-cisterna-explote-con-10-mil-galones-de-combustible" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Bomberos evitan que cami�n cisterna explote con 10 mil galones de combustible</a></h2>
		      	<p class="texto_nota"> (VIDEOS) Los bomberos aplicaron una espuma especial para neutralizar los vapores que emanaba el combustible.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137550/2018/03/21/Bomberos-evitan-que-camion-cisterna-explote-con-10-mil-galones-de-combustible#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137545/2018/03/21/Interiano-asegura-que-ARENA-ha-devuelto-la-esperanza-a-�un-pais-que-estaba-tan-sufrido�"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/TBSO_RFkwNFdmYlhrQUFYaG5aLmpwZw==.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137545/2018/03/21/Interiano-asegura-que-ARENA-ha-devuelto-la-esperanza-a-�un-pais-que-estaba-tan-sufrido�" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Interiano asegura que ARENA ha devuelto la esperanza a �un pa�s que estaba tan sufrido�</a></h2>
		      	<p class="texto_nota"> Expres� que desde la Asamblea Legislativa van a tomar algunas medidas de austeridad y que de hecho ya sus diputados dieron el ejemplo.�</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137545/2018/03/21/Interiano-asegura-que-ARENA-ha-devuelto-la-esperanza-a-�un-pais-que-estaba-tan-sufrido�#comentarios"> (9) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/internacionales/137539/2018/03/21/Se-inmola-el-presunto-autor-de-los-ataques-con-explosivos-en-Texas"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/WVQZ_YXVzdGluLXBhcXVldGVzLWJvbWJhLmpwZWc=.jpeg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/internacionales/137539/2018/03/21/Se-inmola-el-presunto-autor-de-los-ataques-con-explosivos-en-Texas" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Se inmola el presunto autor de los ataques con explosivos en Texas</a></h2>
		      	<p class="texto_nota"> El sospechoso de una oleada de ataques con paquetes bomba que atemorizaron a Austin el mes pasado se inmol&oacute; a primera hora del mi&eacute;rcoles al ser cercado por las autoridades, poniendo fin a un...<a href='http://www.lapagina.com.sv/internacionales/137539/2018/03/21/Se-inmola-el-presunto-autor-de-los-ataques-con-explosivos-en-Texas' style='text-decoration:none;color:#666666;'><i>ampliar</i></a></p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137539/2018/03/21/Se-inmola-el-presunto-autor-de-los-ataques-con-explosivos-en-Texas#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137542/2018/03/21/Ministra-de-Medio-Ambiente-exige-a-los-nuevos-diputados-aprobar-la-Ley-de-Aguas"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/WXDS_RFkwMzRFWldrQUVYOE8tLmpwZw==.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137542/2018/03/21/Ministra-de-Medio-Ambiente-exige-a-los-nuevos-diputados-aprobar-la-Ley-de-Aguas" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Ministra de Medio Ambiente exige a los nuevos diputados aprobar la Ley de Aguas</a></h2>
		      	<p class="texto_nota"> Lina Pohl espera que en la nueva legislatura tomen conciencia que el agua es un recurso fundamental y escaso.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137542/2018/03/21/Ministra-de-Medio-Ambiente-exige-a-los-nuevos-diputados-aprobar-la-Ley-de-Aguas#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/jetset">Jet Set</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/jetset/137549/2018/03/21/Selena-Gomez-recibe-criticas-por-su-cuerpo-y-asi-reacciono"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/GQVP_MzcuanBn.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/jetset/137549/2018/03/21/Selena-Gomez-recibe-criticas-por-su-cuerpo-y-asi-reacciono" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Selena G�mez recibe cr�ticas por su cuerpo y as� reaccion�</a></h2>
		      	<p class="texto_nota"> No es la primera vez que G�mez es v�ctima de este tipo de ataques.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/jetset/137549/2018/03/21/Selena-Gomez-recibe-criticas-por-su-cuerpo-y-asi-reacciono#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/internacionales/137531/2018/03/21/Para-Moscu-el-caso-Skripal-es-un-montaje-de-Londres"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/TFVN_a3JpcGFsLXJlaW5vLXVuaWRvLTY0MHgzNjAuanBn.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/internacionales/137531/2018/03/21/Para-Moscu-el-caso-Skripal-es-un-montaje-de-Londres" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Para Mosc� el caso Skripal es "un montaje de Londres"</a></h2>
		      	<p class="texto_nota"> Las pruebas reales podr�an haber desaparecido ya debido al tiempo que se ha invertido en una ocultaci�n deliberada de los hechos del caso, seg�n la Canciller�a rusa.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137531/2018/03/21/Para-Moscu-el-caso-Skripal-es-un-montaje-de-Londres#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/nacionales/137530/2018/03/21/MARN-pronostica-vientos-para-este-miercoles-"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/AJMH_RFBMRF9ZMnhwYldFdFpXd3RjMkZzZG1Ga2IzSXRO.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/nacionales/137530/2018/03/21/MARN-pronostica-vientos-para-este-miercoles-" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">MARN pronostica vientos para este mi�rcoles </a></h2>
		      	<p class="texto_nota"> Durante el d�a el ambiente estar� c�lido con una temperatura m�xima para San Salvador de 32�C, San Miguel 38� y Santa Ana 34�C.</p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137530/2018/03/21/MARN-pronostica-vientos-para-este-miercoles-#comentarios"> (0) Comentarios</a></div>
		      	<div class='div_puntos'></div>		      	<h1 class="portada"><strong  class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
		      					
	              <a href="http://www.lapagina.com.sv/internacionales/137540/2018/03/21/Se-eleva-la-venta-de-televisores-en-Centroamerica"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/YNJE_U21hcnQtVFYuanBn.jpg" width="340" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>		      	
		      	<h2><a href="http://www.lapagina.com.sv/internacionales/137540/2018/03/21/Se-eleva-la-venta-de-televisores-en-Centroamerica" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Se eleva la venta de televisores en Centroam�rica</a></h2>
		      	<p class="texto_nota"> La venta de televisores en Centroam&eacute;rica increment&oacute; 8% durante los primeros nueve meses de 2017 en comparaci&oacute;n con el mismo periodo de 2016.

Centroam&eacute;rica es un cliente potencial en estos...<a href='http://www.lapagina.com.sv/internacionales/137540/2018/03/21/Se-eleva-la-venta-de-televisores-en-Centroamerica' style='text-decoration:none;color:#666666;'><i>ampliar</i></a></p>
		      	
		      			      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137540/2018/03/21/Se-eleva-la-venta-de-televisores-en-Centroamerica#comentarios"> (0) Comentarios</a></div>
		      	 		     
		    </div>
		    <div id="col_02">
		    					      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/internacionales/137548/2018/03/21/Divulgan-video-con-presunto-intento-de-compra-de-votos-para-Kuczynski"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/LFUU_UEotc2VudGVuY2lhLWEtUFBLLXBvci1kZXVkYS1s.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/internacionales/137548/2018/03/21/Divulgan-video-con-presunto-intento-de-compra-de-votos-para-Kuczynski" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Divulgan video con presunto intento de compra de votos para Kuczynski</a></h2>
				      	

Pedro Pablo Kuczynski (PPK), hizo oficial su renuncia a la Presidencia de la Rep&uacute;blica, luego de que entre ayer y hoy la bancada de Fuerza Popular difundiera un conjunto de audios, en los que se...<a href='http://www.lapagina.com.sv/internacionales/137548/2018/03/21/Divulgan-video-con-presunto-intento-de-compra-de-votos-para-Kuczynski' style='text-decoration:none;color:#666666;'><i>ampliar</i></a>				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137548/2018/03/21/Divulgan-video-con-presunto-intento-de-compra-de-votos-para-Kuczynski#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137543/2018/03/21/�scar-Ortiz-no-buscara-candidatura-presidencial-"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/RJDG_MjMzNUQwQUMtNEY0MS00NkZELTkxOEMtRTFDNzNE.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137543/2018/03/21/�scar-Ortiz-no-buscara-candidatura-presidencial-" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">�scar Ortiz no buscar� candidatura presidencial </a></h2>
				      	El vicepresidente no ha decidido si brindar� su apoyo a la candidatura de Gerson Mart�nez, a quien pidi� hace dos meses que no aceptara el favoritismo y verticalismo de la c�pula.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137543/2018/03/21/�scar-Ortiz-no-buscara-candidatura-presidencial-#comentarios"> (13) Comentarios</a></div>
				      			    			<div class="titulo_notaDestacada"><a  href="http://www.lapagina.com.sv/internacionales" style="color:#ffffff">Internacionales</a></div>
					      <div class="nota_destacada">
						      <h1 class="portada"></h1>
					      					
	              <a href="http://www.lapagina.com.sv/internacionales/137413/2018/03/17/Tigre-se-�come-vivo�-a-su-cuidador-en-un-zoologico-de-China-"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/ZDAH_dGlncmVhdGFjYWN1aWRhZG9yLmpwZw==.jpg" width="253" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>					        
					        <h2><a href="http://www.lapagina.com.sv/internacionales/137413/2018/03/17/Tigre-se-�come-vivo�-a-su-cuidador-en-un-zoologico-de-China-" style="text-decoration:none;color:#ffffff">Tigre se �come vivo� a su cuidador en un zool�gico de China </a></h2>
					        IMAGENES FUERTES.					        <br><br>
					        <div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137413/2018/03/17/Tigre-se-�come-vivo�-a-su-cuidador-en-un-zoologico-de-China-#comentarios">(6) Comentarios</a></div>
					      </div>
		    			<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/internacionales/137547/2018/03/21/Pablo-Kuczynski-renuncia-a-la-presidencia-de-Peru"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/QXQK_UGVkb1BlcnVhc2Rhcy5KUEc=.JPG" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/internacionales/137547/2018/03/21/Pablo-Kuczynski-renuncia-a-la-presidencia-de-Peru" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Pablo Kuczynski renuncia a la presidencia de Per�</a></h2>
				      	La decisi&oacute;n fue tomada luego de una reuni&oacute;n con su gabinete. Ma&ntilde;ana, el Congreso iba a votar su destituci&oacute;n por sus v&iacute;nculos con la constructora brasile&ntilde;a Odebrecht y de comprar votos en el Congreso...<a href='http://www.lapagina.com.sv/internacionales/137547/2018/03/21/Pablo-Kuczynski-renuncia-a-la-presidencia-de-Peru' style='text-decoration:none;color:#666666;'><i>ampliar</i></a>				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137547/2018/03/21/Pablo-Kuczynski-renuncia-a-la-presidencia-de-Peru#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/internacionales/137538/2018/03/21/Cuidador-encuentra-serpiente-con-dos-cabezas-y-dos-corazones"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/YKXK_c2VycGllbnRlZGVkb3NjYWJlemFzLkpQRw==.JPG" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/internacionales/137538/2018/03/21/Cuidador-encuentra-serpiente-con-dos-cabezas-y-dos-corazones" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Cuidador encuentra serpiente con dos cabezas y dos corazones</a></h2>
				      	�VIDEO				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137538/2018/03/21/Cuidador-encuentra-serpiente-con-dos-cabezas-y-dos-corazones#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137551/2018/03/21/Sector-salud-endosa-apoyo-a-Javier-Siman"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/NVPG_bWVkaS5qcGc=.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137551/2018/03/21/Sector-salud-endosa-apoyo-a-Javier-Siman" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Sector salud endosa apoyo a Javier Sim�n</a></h2>
				      	En esta ocasi&oacute;n un grupo de m&eacute;dicos, param&eacute;dicos y enfermeras afines al partido ARENA, dieron apoyo incondicional a Javier Sim&aacute;n, porque creen que es la persona m&aacute;s id&oacute;nea para ocupar la presidencia...<a href='http://www.lapagina.com.sv/nacionales/137551/2018/03/21/Sector-salud-endosa-apoyo-a-Javier-Siman' style='text-decoration:none;color:#666666;'><i>ampliar</i></a>				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137551/2018/03/21/Sector-salud-endosa-apoyo-a-Javier-Siman#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137536/2018/03/21/Obras-en-el-Rancho-Navarra-presentan-un-avance-del-55"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/RTDW_RFlxa29CYldrQVEtSzBYLmpwZw==.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137536/2018/03/21/Obras-en-el-Rancho-Navarra-presentan-un-avance-del-55" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Obras en el Rancho Navarra presentan un avance del 55%</a></h2>
				      	Se tiene previsto que la obra, cuya inversi�n es de m�s de $21 millones,�concluya el pr�ximo mes de abril.�				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137536/2018/03/21/Obras-en-el-Rancho-Navarra-presentan-un-avance-del-55#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137535/2018/03/21/PNC-captura-a-presuntos-traficantes-de-droga-en-la-Tutunichapa"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/JYSM_MGExNWNhNzYtZTA2MS00ZDkxLWFlNGItZDEzNWY3.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137535/2018/03/21/PNC-captura-a-presuntos-traficantes-de-droga-en-la-Tutunichapa" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">PNC captura a presuntos traficantes de droga en la Tutunichapa</a></h2>
				      	En otro procedimiento, personal de Investigaciones captur� a Henry Adiel D�az Corado por simulaci�n de delito.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137535/2018/03/21/PNC-captura-a-presuntos-traficantes-de-droga-en-la-Tutunichapa#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137534/2018/03/21/Al-menos-diez-pandilleros-detenidos-por-el-delito-de-homicidio"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/FBUF_Q2FwdHVyYXNhc2RhczIzMy5KUEc=.JPG" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137534/2018/03/21/Al-menos-diez-pandilleros-detenidos-por-el-delito-de-homicidio" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Al menos diez pandilleros detenidos por el delito de homicidio</a></h2>
				      	La PNC realiz� diez capturas de miembros de pandillas y la FGR orden� la captura de 31 sujetos pertenecientes a estructuras criminales.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137534/2018/03/21/Al-menos-diez-pandilleros-detenidos-por-el-delito-de-homicidio#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/deportes">Deportes</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/deportes/137533/2018/03/21/Xavi-Alonso-podria-ir-a-la-carcel"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/TQWR_MTQ3NjcwOTA2Ml8wNjYwNzhfMTQ3NjcxNDA5NV9u.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/deportes/137533/2018/03/21/Xavi-Alonso-podria-ir-a-la-carcel" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Xavi Alonso podr�a ir a la c�rcel</a></h2>
				      	Entre 2009 y 2012, Alonso, seg�n la Fiscal�a, explot� su imagen a distintas empresas que le contrataban con la ayuda de otros dos acusados sin hacer &ldquo;uso real&rdquo; de la sociedad.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/deportes/137533/2018/03/21/Xavi-Alonso-podria-ir-a-la-carcel#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/nacionales">Nacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/nacionales/137541/2018/03/21/Raul-Mijango-Esto-es-parte-de-un-show-politico-de-la-Fiscalia"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/TJCT_TWlqYW5nb2FzZGFzZC5KUEc=.JPG" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/nacionales/137541/2018/03/21/Raul-Mijango-Esto-es-parte-de-un-show-politico-de-la-Fiscalia" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Ra�l Mijango: "Esto es parte de un show pol�tico de la Fiscal�a"</a></h2>
				      	La reacci�n de Mijango se da en el marco de que la C�mara Especializada de lo Penal anul� el juicio que se llev� a cabo contra los procesados por la tregua de pandillas.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/nacionales/137541/2018/03/21/Raul-Mijango-Esto-es-parte-de-un-show-politico-de-la-Fiscalia#comentarios"> (0) Comentarios</a></div>
				      	<div class='div_puntos'></div>				      	<h1 class="portada"><strong class="seccion"><a href="http://www.lapagina.com.sv/internacionales">Internacionales</a></strong>  </h1>
				      					
	              <a href="http://www.lapagina.com.sv/internacionales/137528/2018/03/21/Papa-Francisco-admite-renuncia-del-prefecto-de-comunicaciones-tras-polemica-por-carta-de-Benedicto-XVI"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/ARPK_OWE0OWJhYzJlMzAxZGEzN2Q3NmFlMWM4ZDE1ZDNh.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>				      	
				      	<h2><a href="http://www.lapagina.com.sv/internacionales/137528/2018/03/21/Papa-Francisco-admite-renuncia-del-prefecto-de-comunicaciones-tras-polemica-por-carta-de-Benedicto-XVI" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Papa Francisco admite renuncia del prefecto de comunicaciones, tras pol�mica por carta de Benedicto XVI</a></h2>
				      	No obstante, monse�or Vigan� permanecer� en el Dicasterio como asesor del nuevo prefecto.				      	<br><br>
				      					      	<div class="boton_verComentarios"><a href="http://www.lapagina.com.sv/internacionales/137528/2018/03/21/Papa-Francisco-admite-renuncia-del-prefecto-de-comunicaciones-tras-polemica-por-carta-de-Benedicto-XVI#comentarios"> (0) Comentarios</a></div>
				      			    </div>
		  </div>
		<div id="col_derecha" >
<!---	<div class="especial_ld">
			<a href="https://goo.gl/tBZLdc" target="_blank"><img src="http://www.lapagina.com.sv/campo_pagado/comunicado_15022018.jpg" border="0"></a>
			
		</div> 
 
	<div class="div_puntos"></div>  
	
	<div class="especial_campain">
			<div class="tituloesp">
				<p class="tes"> #HacemosMasPorLaGente </p>
			</div>
			<iframe width="290" height="163" src="https://www.youtube-nocookie.com/embed/ivq9vdHBnpI?rel=0&amp;showinfo=0" frameborder="0" allow="autoplay; encrypted-media" allowfullscreen></iframe>
			
		</div> 
 
	<div class="div_puntos"></div>  
<!---	<div class="especial_ld">
			<a href="https://goo.gl/tm6Wxn" target="_blank"><img src="http://www.lapagina.com.sv/campo_pagado/comunicado_15022018.jpg" border="0"></a>
			
		</div> 
 
	<div class="div_puntos"></div> ---> 
	 
    				
	              <a href="http://www.lapagina.com.sv/internacionales/137537/2018/03/21/Dama-de-compania-filtro-video-de-su-asesino"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/LRHM_ZXNwZXJhbWUtdW4tcG9xdWl0by1hc2ktcHVlZG8t.jpg" width="300" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>            <h2><a href="http://www.lapagina.com.sv/internacionales/137537/2018/03/21/Dama-de-compania-filtro-video-de-su-asesino" style="text-decoration:none;color:#8E151F;font-size:px;line-height:px">Dama de compa��a filtr� video de su asesino</a></h2>
    Con golpes y signos de tortura, fue encontrado el cuerpo de Kenni el pasado 25 de febrero. Su cad&aacute;ver fue hallado tirado en una calle, frente a una escuela. En su rostro le echaron &aacute;cido, luego le...<a href='http://www.lapagina.com.sv/internacionales/137537/2018/03/21/Dama-de-compania-filtro-video-de-su-asesino' style='text-decoration:none;color:#666666;'><i>ampliar</i></a>            <br><br>
            <div class="boton_verComentarios">
                <a href="http://www.lapagina.com.sv/internacionales/137537/2018/03/21/Dama-de-compania-filtro-video-de-su-asesino#comentarios">(0) Comentarios</a>
            </div>
            <div class="div_puntos"></div>
        
    <!-- Script DOUBLECLICK - Banner_lateral_izquierdo_1-->
    <!-- lateral_derecho_1 -->
    
    <script type='text/javascript'>
        GA_googleFillSlot("lateral_derecho_1");
    </script>
    <!-- Fin Script DOUBLECLICK - Banner_lateral_izquierdo_1-->

     
    <div class="wsbotton"> 
                  
	<div class="div_puntos"></div>

                            <div id="rotador_0" style="display:none">
                            <p class="titulosSecciones"><a href="http://www.lapagina.com.sv/cultura" style="color:#ffffff">Cultura</a></p>
                            <div class="contenedor_ocio">
	                             <p class="copete"></p>
                            <div class="img_rota"> 				
	              <a href="http://www.lapagina.com.sv/cultura/137378/2018/03/16/Hombre-viaja-por-Mexico-curando-a-perros-callejeros--"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/FBXW_ZmFjZWJvb2stcGVycm9zMi0xNTIwNzkxMDM0Lmpw.jpg" width="276" style="margin-bottom:0px;margin-right:5px;" alt=""/></a> 
		                        </div>
	                            <div class="titular_rota"><h2 class="ocio"><a href="http://www.lapagina.com.sv/cultura/137378/2018/03/16/Hombre-viaja-por-Mexico-curando-a-perros-callejeros--" style="text-decoration:none;color:#555555">Hombre viaja por M�xico curando a perros callejeros  </a></h2>
	                            </div>
		                         <p class="font12">VIDEO VIRAL.</p>              
            				</div>
        				</div>
                            <div id="rotador_1" style="display:none">
                            <p class="titulosSecciones"><a href="http://www.lapagina.com.sv/jetset" style="color:#ffffff">Jet Set</a></p>
                            <div class="contenedor_ocio">
	                             <p class="copete"></p>
                            <div class="img_rota"> 				
	              <a href="http://www.lapagina.com.sv/jetset/137349/2018/03/15/Coqueteo-con-una-sexy-modelo-su-novia-lo-descubrio-y-lo-dejo-expuesto--"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/IAET_NzUyMTQuanBn.jpg" width="276" style="margin-bottom:0px;margin-right:5px;" alt=""/></a> 
		                        </div>
	                            <div class="titular_rota"><h2 class="ocio"><a href="http://www.lapagina.com.sv/jetset/137349/2018/03/15/Coqueteo-con-una-sexy-modelo-su-novia-lo-descubrio-y-lo-dejo-expuesto--" style="text-decoration:none;color:#555555">Coquete� con una sexy modelo, su novia lo descubri� y lo dej� expuesto  </a></h2>
	                            </div>
		                         <p class="font12">El joven respondi&oacute; con un p&iacute;caro mensaje a una publicaci&oacute;n de la argentina...<a href='http://www.lapagina.com.sv/jetset/137349/2018/03/15/Coqueteo-con-una-sexy-modelo-su-novia-lo-descubrio-y-lo-dejo-expuesto--' style='text-decoration:none;color:#666666;'><i>ampliar</i></a></p>              
            				</div>
        				</div>
                            <div id="rotador_2" style="display:none">
                            <p class="titulosSecciones"><a href="http://www.lapagina.com.sv/curiosidades" style="color:#ffffff">Curiosidades</a></p>
                            <div class="contenedor_ocio">
	                             <p class="copete">COLOMBIA</p>
                            <div class="img_rota"> 				
	              <a href="http://www.lapagina.com.sv/curiosidades/137348/2018/03/15/Motorista-atrapa-a-ladron-con-las-puertas-del-bus-"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/FOFA_bGFkcm9uYnVzLnBuZw==.png" width="276" style="margin-bottom:0px;margin-right:5px;" alt=""/></a> 
		                        </div>
	                            <div class="titular_rota"><h2 class="ocio"><a href="http://www.lapagina.com.sv/curiosidades/137348/2018/03/15/Motorista-atrapa-a-ladron-con-las-puertas-del-bus-" style="text-decoration:none;color:#555555">Motorista atrapa a ladr�n con las puertas del bus </a></h2>
	                            </div>
		                         <p class="font12">�VIDEO</p>              
            				</div>
        				</div>
                            <div class="botones_ocio"><a href="javascript:rotar(0);">&lt;    &nbsp;ANTERIOR</a>&nbsp;  |&nbsp; <a href="javascript:rotar(1);">SIGUIENTE&nbsp;    &gt;</a></div>
                        <script>
                              			document.getElementById("rotador_0").style.display="inline";
                              			var actual = 0;
                              			function rotar(sentido){
                              				ant = actual;
                              				if (sentido==0){
                              					if (actual==0) actual = 2;
                              					else actual--;
                              				}
                              				else if (actual==2) actual = 0;
                              					 else actual++;
                              				document.getElementById("rotador_"+ant).style.display="none";
                              				document.getElementById("rotador_"+actual).style.display="inline";
                              			}
                        </script>
</div>

<div class="div_puntos"></div>

    <!-- lateral_derecho_4 -->
    <script type='text/javascript'>
        GA_googleFillSlot("lateral_derecho_4");
    </script>

<div class="div_puntos"></div>

	<!--
  SELECT n.id, n.titular, n.galeria, n.fecha_modificacion, s.nombre
  FROM lomas l, noticias n
  JOIN secciones s ON n.seccion = s.id
  WHERE n.id = l.id_noticia
    AND l.tipo = 'leido'
  ORDER BY l.orden ASC--><script>
	function ver_lomas(n){
		if (n==0){
			document.getElementById("lomascomentado").style.display="none";
			document.getElementById("lomasleido").style.display="inline";
			document.getElementById("pes0b").style.display="none";
			document.getElementById("pes1b").style.display="none";
			document.getElementById("pes0a").style.display="inline";
			document.getElementById("pes1a").style.display="inline";
		}
		else{
			document.getElementById("lomascomentado").style.display="inline";
			document.getElementById("lomasleido").style.display="none";
			document.getElementById("pes0a").style.display="none";
			document.getElementById("pes1a").style.display="none";
			document.getElementById("pes0b").style.display="inline";
			document.getElementById("pes1b").style.display="inline";
		}
	}
</script>
<div id="lomas">
<div id="pes1a" class="pestanias_select" style="cursor:pointer;float:left" onclick="ver_lomas(0);">
	<table width="110" border="0" cellpadding="0" cellspacing="0" class="pestaniaSelect">
	    <tr>
	      <td width="7"><img src="http://www.lapagina.com.sv/images/pestanias/on_izq.gif" width="7" height="28" /></td>
	      <td background="http://www.lapagina.com.sv/images/pestanias/on_back.gif"><div align="center">LO M&Aacute;S LE&Iacute;DO </div></td>
	      <td width="9"><img src="http://www.lapagina.com.sv/images/pestanias/on_der.gif" width="9" height="28" /></td>
	    </tr>
	</table>
</div>
<div id="pes0a" class="pestanias" style="cursor:pointer;" onclick="ver_lomas(1);">
<table width="140" border="0" cellpadding="0" cellspacing="0" class="pestaniaNoSelect">
	            <tr>
	              <td width="7"><img src="http://www.lapagina.com.sv/images/pestanias/off_izq.gif" width="7" height="28" /></td>
	              <td background="http://www.lapagina.com.sv/images/pestanias/off_back.gif"><div align="center">LO M&Aacute;S COMENTADO </div></td>
	              <td width="9"><img src="http://www.lapagina.com.sv/images/pestanias/off_der.gif" width="9" height="28" /></td>
	            </tr>
	        </table>
</div>
<div id="pes1b" class="pestanias_select" style="cursor:pointer;float:left;display:none" onclick="ver_lomas(0);">
	<table width="110" border="0" cellpadding="0" cellspacing="0" class="pestaniaNoSelect">
        <tr>
          <td width="7"><img src="http://www.lapagina.com.sv/images/pestanias/off_izq.gif" width="7" height="28" /></td>
          <td background="http://www.lapagina.com.sv/images/pestanias/off_back.gif"><div align="center">LO M&Aacute;S LE&Iacute;DO </div></td>
          <td width="9"><img src="http://www.lapagina.com.sv/images/pestanias/off_der.gif" width="9" height="28" /></td>
        </tr>
    </table>
</div>
<div id="pes0b" class="pestanias" style="cursor:pointer;display:none;" onclick="ver_lomas(1);">
	<table width="140" border="0" cellpadding="0" cellspacing="0" class="pestaniaSelect">
	    <tr>
	      <td width="7"><img src="http://www.lapagina.com.sv/images/pestanias/on_izq.gif" width="7" height="28" /></td>
	      <td background="http://www.lapagina.com.sv/images/pestanias/on_back.gif"><div align="center">Lo m&Aacute;s comentado </div></td>
	      <td width="9"><img src="http://www.lapagina.com.sv/images/pestanias/on_der.gif" width="9" height="28" /></td>
	    </tr>
	</table>
</div>

	<div id="lomasleido" style="display:inline">
  	  	  <a href="http://www.lapagina.com.sv/jetset/136794/2018/02/23/Filtran-video-erotico-de-sexy-candidata-a-alcaldesa-" style="text-decoration:none">
  	  	<div class="lineas_contenidos"  style="cursor:pointer;">
  	  		<p class="lomasClaro">Filtran video er�tico de sexy "candidata" a alcaldesa </p>
  	  	</div>
  	  </a>
  	
  		  <a href="http://www.lapagina.com.sv/nacionales/136931/2018/02/28/Camaras-del-Hospital-San-Rafael-captan-actividad-paranormal-frente-a-la-morgue" style="color:#999999;text-decoration:none">
		  
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">C�maras del Hospital San Rafael captan actividad paranormal frente a la morgue</p>
	  	</div>
	  </a>
	
		  <a href="http://www.lapagina.com.sv/internacionales/136793/2018/02/23/Trump-reclama-a-El-Salvador-por-tomar-su-dinero" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">
	  			Trump reclama a El Salvador por "tomar su dinero"	  		</p>
	  	</div>
	  </a>
		  <a href="http://www.lapagina.com.sv/nacionales/136817/2018/02/24/Gobierno-de-El-Salvador-condena-declaraciones-de-Donald-Trump" style="color:#999999;text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">Gobierno de El Salvador condena declaraciones de Donald Trump</p>
	  	</div>
	  </a>
	
		  <a href="http://www.lapagina.com.sv/nacionales/136915/2018/02/27/Capturan-a-subinspector-de-la-PNC-por-muerte-de-su-esposa" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">Capturan a subinspector de la PNC por muerte de su esposa</p>
	  	</div>
	  </a>
		  <a href="http://www.lapagina.com.sv/nacionales/136857/2018/02/26/PNC-cree-haber-encontrado-tumba-donde-estaria-el-cuerpo-de-la-agente-Carla-Ayala" style="color:#999999;text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">PNC cree haber encontrado tumba donde estar�a el cuerpo de la agente Carla Ayala</p>
	  	</div>
	  </a>
		  <a href="http://www.lapagina.com.sv/internacionales/136923/2018/02/28/Trump-solo-bajo-un-gran-paraguas-y-deja-a-su-mujer-e-hijo-expuestos-a-la-lluvia" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">Trump solo bajo un gran paraguas y deja a su mujer e hijo expuestos a la lluvia</p>
	  	</div>
	  </a>
	
  </div>
  <div id="lomascomentado" style="display:none">
  		  <a href="http://www.lapagina.com.sv/internacionales/136793/2018/02/23/Trump-reclama-a-El-Salvador-por-tomar-su-dinero" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">Trump reclama a El Salvador por "tomar su dinero"</p>
	  	</div>
	  </a>
		  <a href="http://www.lapagina.com.sv/nacionales/136810/2018/02/23/Alta-funcionaria-de-Trump-hara-gira-por-Triangulo-Norte-menos-por-El-Salvador" style="color:#999999;text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">Alta funcionaria de Trump har� gira por Tri�ngulo Norte, menos por El Salvador</p>
	  	</div>
	  </a>
	  
		  <a href="http://www.lapagina.com.sv/nacionales/136817/2018/02/24/Gobierno-de-El-Salvador-condena-declaraciones-de-Donald-Trump" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">Gobierno de El Salvador condena declaraciones de Donald Trump</p>
	  	</div>
	  </a>
	  	  <a href="http://www.lapagina.com.sv/nacionales/136931/2018/02/28/Camaras-del-Hospital-San-Rafael-captan-actividad-paranormal-frente-a-la-morgue" style="color:#999999;text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">C�maras del Hospital San Rafael captan actividad paranormal frente a la morgue</p>
	  	</div>
	  </a>
	  
		  <a href="http://www.lapagina.com.sv/nacionales/136927/2018/02/28/Por-que-le-tienen-miedo-a-Jose-Luis-Merino-se-cuestiona-candidato-del-FMLN" style="text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasClaro">"�Por qu� le tienen miedo a Jos� Luis Merino?", se cuestiona candidato del FMLN</p>
	  	</div>
	  </a>
	  	  <a href="http://www.lapagina.com.sv/nacionales/136913/2018/02/27/PNC-vuelve-a-perder-el-rastro-de-Carla-Ayala-Cuerpo-exhumado-es-de-una-mujer-que-murio-a-los-91-anos" style="color:#999999;text-decoration:none">
	  	<div class="lineas_contenidos" style="cursor:pointer;">
	  		<p class="lomasOscuro">PNC vuelve a perder el rastro de Carla Ayala: Cuerpo exhumado es de una mujer que muri� a los 91 a�os</p>
	  	</div>
	  </a>
	  
		  <a href="http://www.lapagina.com.sv/nacionales/136895/2018/02/27/Maria-Isabel-Rodriguez-se-pronuncia-en-contra-del-voto-nulo" style="text-decoration:none"><div class="lineas_contenidos" style="cursor:pointer;">Mar�a Isabel Rodr�guez se pronuncia en contra del voto nulo</div></a>
	  		</td>
	  	</tr>
	  </table>
  </div>
</div>

	
		
		<div class="div_puntos"></div>
        
        <script type='text/javascript'>
            GA_googleFillSlot("lateral_derecho_2");
        </script>
        
        <script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>

<div class="div_puntos"></div>

    <p class="titulosSecciones">
        <a href="http://www.lapagina.com.sv/entrevistas" style="color:#ffffff">
  		LA ENTREVISTA
        </a>
    </p>
        <div class="contenedor_entrevistas">
        				
	              <a href="http://www.lapagina.com.sv/entrevistas/137527/Salvadorena-representa-al-pais-en-evento-cientifico-mundial-en-EEUU"><img class="portada" src="http://www.lapagina.com.sv/userfiles/Mar_2018/UMYU_RXZlbHluVVNBLmpwZw==.jpg" width="270" style="margin-bottom:0px;margin-right:5px;" alt=""/></a>        <p class="copete"></p>
        <h2><a href="http://www.lapagina.com.sv/entrevistas/137527/Salvadorena-representa-al-pais-en-evento-cientifico-mundial-en-EEUU" style="text-decoration:none;color:#555555">Salvadore�a representa al pa�s en evento cient�fico mundial en EE.UU</a></h2>
        Una joven salvadore&ntilde;a, originaria de Ciudad Delgado representa a la Universidad de Illinois, Estados Unidos y a El Salvador en el Global Food Security Symposium 2018, un evento mundial, en el que se...<a href='http://www.lapagina.com.sv/entrevistas/137527/Salvadorena-representa-al-pais-en-evento-cientifico-mundial-en-EEUU' style='text-decoration:none;color:#666666;'><i>ampliar</i></a>        </div>

<div class="div_puntos"></div>

            <!-- lateral_derecho_3 -->
            <script type='text/javascript'>
                GA_googleFillSlot("lateral_derecho_3");
            </script>        

<div class="div_puntos"></div>
        <p class="titulosSecciones">OPINION</p>
                    <div class="opinion">
                    <table width="302" border="0" cellspacing="4" cellpadding="0" class="">
                        <tr valign="top">
                            <td width="48">
                                <img src="http://www.lapagina.com.sv/userfiles/autores/NPUW_U1ZDWl9jMlZ1YjNJdWFuQmwuanBl.jpe" width="70" height="70" class="img_marcoGrisOscuro" />
                            </td>
                            <td>
                                <p class="titulo"><a href="http://www.lapagina.com.sv/editoriales/137532/Esta-derrotado-el-FMLN" style="text-decoration:none;color:#555555">�Est� derrotado el FMLN?</a></p>
                                <p class="nombre">Carlos Argueta</p>
                            </td>
                        </tr>
                    </table>
                </div>
                    <div class="opinion">
                    <table width="302" border="0" cellspacing="4" cellpadding="0" class="tablaOscura">
                        <tr valign="top">
                            <td width="48">
                                <img src="http://www.lapagina.com.sv/userfiles/autores/NPUW_U1ZDWl9jMlZ1YjNJdWFuQmwuanBl.jpe" width="70" height="70" class="img_marcoGrisOscuro" />
                            </td>
                            <td>
                                <p class="titulo"><a href="http://www.lapagina.com.sv/editoriales/137256/No-fue-la-corrupcion-ni-lo-economico-Es-la-falta-de-alianzas-" style="text-decoration:none;color:#555555">No fue la corrupci�n, ni lo econ�mico. Es la falta de alianzas </a></p>
                                <p class="nombre">Carlos Argueta</p>
                            </td>
                        </tr>
                    </table>
                </div>
                    <div class="opinion">
                    <table width="302" border="0" cellspacing="4" cellpadding="0" class="">
                        <tr valign="top">
                            <td width="48">
                                <img src="http://www.lapagina.com.sv/userfiles/autores/OFCH_Rk9UT19EUi5fRkpGLkpQRw==.JPG" width="70" height="70" class="img_marcoGrisOscuro" />
                            </td>
                            <td>
                                <p class="titulo"><a href="http://www.lapagina.com.sv/editoriales/137262/El-Salvador-no-es-laboratorio-de-los-populismos" style="text-decoration:none;color:#555555">El Salvador no es laboratorio de los populismos</a></p>
                                <p class="nombre">Francisco Jos� Ferm�n </p>
                            </td>
                        </tr>
                    </table>
                </div>
                    <div class="opinion">
                    <table width="302" border="0" cellspacing="4" cellpadding="0" class="tablaOscura">
                        <tr valign="top">
                            <td width="48">
                                <img src="http://www.lapagina.com.sv/userfiles/autores/OFCH_Rk9UT19EUi5fRkpGLkpQRw==.JPG" width="70" height="70" class="img_marcoGrisOscuro" />
                            </td>
                            <td>
                                <p class="titulo"><a href="http://www.lapagina.com.sv/editoriales/137167/El-poder-soberano-se-manifiesta-" style="text-decoration:none;color:#555555">El poder soberano se manifiesta </a></p>
                                <p class="nombre">Francisco Jos� Ferm�n </p>
                            </td>
                        </tr>
                    </table>
                </div>
                <div class="contenedor_botones">
                <p class="boton"><a href="http://www.lapagina.com.sv/opinion">VER TODAS</a></p>
            </div>


           
<div class="div_puntos"></div>
 
    <!-- lateral_derecho_5 -->
    <div>
    <script type='text/javascript'>
        GA_googleFillSlot("lateral_derecho_5");
    </script>            
    </div>
<div class="div_puntos"></div>
<div class="encuesta" data-sticky_column>
    <script>
	var votado_inc = 0;
	function enviar_votacion(){
		if (votado_inc) alert("Ya ha votado, gracias por participar");
		else {
			seleccion = false;
			for (i=0;i<document.getElementById("encuesta_inc").resp.length;i++) 
				if (document.getElementById("encuesta_inc").resp[i].checked) seleccion = true;
			if (seleccion)	document.getElementById("encuesta_inc").submit();
			else alert("Seleccione una respuesta.");
		}		
	}
</script>

<div class="encuentas">
	<p class="titulosSecciones">ENCUESTA</p>
	<div class="top_encuesta">
      <h4>�Cree que el m�todo de conteo de votos desarrollado por el TSE es transparente y leg�timo? </h4>
  	</div>
  		<form id="encuesta_inc" method="POST" target="" action="http://www.lapagina.com.sv/res_encuesta.php?id_encuesta=747">
  		  	<div class="respuestas">
	  	<label>
	  		<input type="radio" name="resp" id="resp1" value="1" />
	  		<i></i>
	  		<span class="respuesta"><label for="resp1">No me interesa</label></span>
  	</div>
  	<div class="respuestas">
	  	<label>
	  		<input type="radio" name="resp" id="resp2" value="2" />
	  		<i></i>
	  		<span class="respuesta"><label for="resp2">Si lo es</label></span>
  	</div>
  	<div class="respuestas">
	  	<label>
	  		<input type="radio" name="resp" id="resp3" value="3" />
	  		<i></i>
	  		<span class="respuesta"><label for="resp3">Por supuesto que no </label></span>
  	</div>
<div class="encuesta_boton">
	<a class="encuesta" href="javascript:enviar_votacion()">VOTAR</a>
</div>
  </form>
  <div class="resultados">
      <p class="boton"><a href="http://www.lapagina.com.sv/res_encuesta.php?id_encuesta=747">Ver resultados</a></p>
</div>
</div>
</div>
<div class="div_puntos"></div>

<iframe src="https://www.facebook.com/plugins/page.php?href=https%3A%2F%2Fwww.facebook.com%2FDiarioLaPaginaSV%2F&tabs=timeline&width=300&height=600&small_header=true&adapt_container_width=true&hide_cover=false&show_facepile=false&appId=305661439786665" width="300" height="600" style="border:none;overflow:hidden" scrolling="no" frameborder="0" allowTransparency="true"></iframe>

<div class="div_puntos"></div>
    </div>
		  <div class="end"></div>
		</div>

<div id="base_anuncios_google">
        <!-- Banners cintillos -->
    <div id="bannerPequeno">
        <div class="bannerPeq">
            <!-- footer_cintillo_izquierda -->
            <script type='text/javascript'>
                GA_googleFillSlot("footer_Izq");
            </script>
        </div>

        <div class="bannerPeq">
            <!-- footer_cintillo_central -->
            <script type='text/javascript'>
                GA_googleFillSlot("footer_centro");
            </script>
        </div>

        <div class="bannerPeq">
            <!-- footer_cintillo_derecha -->
            <script type='text/javascript'>
                GA_googleFillSlot("footer_derecha");
            </script>
        </div>

        <div class="end"></div>
    </div>
</div>
<div id="base_recomendamos">
</div>
<div class="base_menu">
  <div id="menu_bottom">
    <p class="botones"><a href="http://www.lapagina.com.sv/portada"  style='color:#ffffff'>PORTADA</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/nacionales" >NACIONALES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/internacionales" >INTERNACIONALES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/entrevistas" >entrevistas</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/empresarial" >empresarial</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/opinion" >OPINI&Oacute;N</a> </p>
    <p class="botones"><a href="http://www.lapagina.com.sv/cultura" >CULTURA</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/deportes" >DEPORTES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/jetset" >JET SET</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/curiosidades"  ?>Curiosidades</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/editoriales">EDITORIALES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/boletines.php">BOLETINES</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/rss.php">RSS</a></p>
    <p class="botones"><a href="http://www.lapagina.com.sv/hemeroteca.php">HEMEROTECA</a></p>
    
  
  </div>
</div><footer>
<div id="base_footer">
  <div id="footer">
    <table width="995" border="0" cellpadding="0" cellspacing="0">
      <tr>
        <td width="260"><a href="http://www.lapagina.com.sv/"portada"><img src="http://www.lapagina.com.sv/images/footer/logopie-1.png" width="260" height="71" border="0" /></a></td>
        <td>TODOS LOS DERECHOS RESERVADOS   
      </td>
        <td width="203"><a href="#"><img src="http://www.lapagina.com.sv/images/footer/Grupo_footer.png" width="203" height="71" border="0" /></a></td>
      </tr>
    </table>
  </div>
</div>
<div class="base_menu">
  <div id="menu_bottom">
    <p class="botones" style="font-size:8pt; text-transform:none; font-weight:normal"><b>Diario La P&aacute;gina</b>. Direcci&oacute;n: Calle La Ceiba 272, Colonia Escalon, San Salvador, El Salvador. Tel&eacute;fono: (503) 2243-8969 | (503) 2246-0616 - Cont&aacute;ctenos a <a href="mailto:redaccion@lapagina.com.sv">redaccion@lapagina.com.sv</a></p>
  </div>
</div>
<!-- Quantcast Tag -->
<script type="text/javascript">
var _qevents = _qevents || [];

(function() {
var elem = document.createElement('script');
elem.src = (document.location.protocol == "https:" ? "https://secure" : "http://edge") + ".quantserve.com/quant.js";
elem.async = true;
elem.type = "text/javascript";
var scpt = document.getElementsByTagName('script')[0];
scpt.parentNode.insertBefore(elem, scpt);
})();

_qevents.push({
qacct:"p-KLe-tShcVVh20"
});
</script>

<noscript>
<div style="display:none;">
<img src="//pixel.quantserve.com/pixel/p-KLe-tShcVVh20.gif" border="0" height="1" width="1" alt="Quantcast"/>
</div>
</noscript>
<!-- End Quantcast tag -->
</footer>


</body>
</html>