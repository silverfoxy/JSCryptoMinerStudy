<!DOCTYPE html>
<!--[if lt IE 7]>      <html class="no-js lt-ie9 lt-ie8 lt-ie7"> <![endif]-->
<!--[if IE 7]>         <html class="no-js lt-ie9 lt-ie8"> <![endif]-->
<!--[if IE 8]>         <html class="no-js lt-ie9"> <![endif]-->
<!--[if gt IE 8]><!-->
<html class="no-js">
<!--<![endif]-->
<head>
<meta charset="utf-8">
<meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
<title>El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal! | Canal 12</title>
<meta name="viewport" content="width=device-width, initial-scale=1">
<!-- Google / Inicio -->
<meta name="description" content="Noticias de El Salvador y el mundo, tenemos las últimas noticias sobre actualidad, deportes, entretenimiento y mucho más en Canal 3.">
<meta name="keywords" content="Noticias de El Salvador, actualidad, deportes, entretenimiento"/>
<meta name="news_keywords" content="Noticias de El Salvador, actualidad, deportes, entretenimiento"/>
<meta name="language" content="es" />
<meta name="robots" content="index,follow"/>
<meta name="googlebot" content="index, follow" />
<meta name="organization" content="Red El Salvador S.A." />
<meta name="revisit-after" content="1 day" />
<meta name="author" content="Canal 12" />
<meta name="copyright" content="©2015 www.canal12.com.sv" />
<meta name="origen" content='Canal 12' />
<meta name="locality" content="San Salvador, El Salvador" />
<meta name="distribution" content="global" />
<link rel="image_src" href="http://cdn.canal12.com.sv/sites/common/img/logo_canal12.png" />
<meta name="dcterms.abstract" content="El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal! - Noticias de El Salvador y el mundo, tenemos las últimas noticias sobre actualidad, deportes, entretenimiento y mucho más en Canal 3." />
<meta name="dcterms.rightsHolder" content="Canal 12">
<link rel="canonical" href="http://canal12.com.sv/"/>
<!-- Google / Fin -->
<!-- Open Graph / Inicio -->
<meta property="og:title" content="El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal! - Canal 12"/>
<meta property="og:site_name" content="Canal 12"/>
<meta property="og:url" content="http://canal12.com.sv/"/>
<meta property="og:description" content="Noticias de El Salvador y el mundo, tenemos las últimas noticias sobre actualidad, deportes, entretenimiento y mucho más en Canal 3."/>
<meta property="og:image" content="http://cdn.canal12.com.sv/sites/common/img/logo_canal12.png"/>
<meta property="fb:app_id" content="263691693659158"/>
<meta property="og:type" content="website"/>
<meta property="article:author" content="https://www.facebook.com/CanalDoceSV" />
<meta property="article:publisher" content="https://www.facebook.com/CanalDoceSV" />
<meta property="article:modified_time" content="2018-03-21 07:03:58 -06:00"/>
<meta property="article:section" content="El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal!"/>
<!-- Open Graph / Fin -->
<!-- Twitter Card / Inicio -->
<meta name="twitter:site" content="@Canal_12" />
<meta name="twitter:title" content="El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal! - Canal 12"/>
<meta name="twitter:description" content="El Salvador en vivo ¡Disfruta lo mejor de nuestra programación y conéctate a nuestra señal! - Noticias de El Salvador y el mundo, tenemos las últimas noticias sobre actualidad, deportes, entretenimiento y mucho más en Canal 3." />
<meta name="twitter:creator" content="@Canal_12">
<meta name="twitter:domain" content="canal12.com.sv">
<meta name="twitter:card" content="summary_large_image"/>
<meta name="twitter:image" content="http://cdn.canal12.com.sv/sites/common/img/logo_canal12.png"/>
<!-- Twitter Card / Fin -->
<link rel="shortcut icon" href="/favicon.ico">
<link rel="apple-touch-icon" sizes="57x57" href="/apple-touch-icon-57x57.png">
<link rel="apple-touch-icon" sizes="60x60" href="/apple-touch-icon-60x60.png">
<link rel="apple-touch-icon" sizes="72x72" href="/apple-touch-icon-72x72.png">
<link rel="apple-touch-icon" sizes="76x76" href="/apple-touch-icon-76x76.png">
<link rel="apple-touch-icon" sizes="114x114" href="/apple-touch-icon-114x114.png">
<link rel="apple-touch-icon" sizes="120x120" href="/apple-touch-icon-120x120.png">
<link rel="apple-touch-icon" sizes="144x144" href="/apple-touch-icon-144x144.png">
<link rel="apple-touch-icon" sizes="152x152" href="/apple-touch-icon-152x152.png">
<link rel="apple-touch-icon" sizes="180x180" href="/apple-touch-icon-180x180.png">
<link rel="icon" type="image/png" href="/favicon-32x32.png" sizes="32x32">
<link rel="icon" type="image/png" href="/favicon-194x194.png" sizes="194x194">
<link rel="icon" type="image/png" href="/favicon-96x96.png" sizes="96x96">
<link rel="icon" type="image/png" href="/android-chrome-192x192.png" sizes="192x192">
<link rel="icon" type="image/png" href="/favicon-16x16.png" sizes="16x16">
<link rel="manifest" href="/manifest.json">
<link rel="mask-icon" href="/safari-pinned-tab.svg" color="#2d89ef">
<meta name="msapplication-TileColor" content="#2d89ef">
<meta name="msapplication-TileImage" content="/mstile-144x144.png">
<meta name="theme-color" content="#6cbced">
<link rel="stylesheet" href="http://cdn.canal12.com.sv/sites/common/css/bootstrap.min.css">
<link rel="stylesheet" href="http://cdn.canal12.com.sv/sites/common/css/default.css">
<link rel="stylesheet" href="http://cdn.canal12.com.sv/sites/common/css/jquery.mobile-1.4.5.min.css">
<link rel="stylesheet" href="http://cdn.canal12.com.sv/sites/canal9/css/default.css">
<script src="http://cdn.canal12.com.sv/sites/common/js/vendor/jquery-1.11.0.min.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/vendor/jquery.mobile.custom.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/vendor/bootstrap.min.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/vendor/modernizr-2.6.2.min.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/vendor/swfobject.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/jquery.lazyload.js"></script>
<script src="http://cdn.canal12.com.sv/sites/common/js/default.js"></script>
<script src="http://cdn.canal12.com.sv/sites/canal9/js/home_principal.js"></script>

<!--
<script src="http://aklc.img.e-planning.net/layers/hbdfp.js" id="hbepl" async="" data-isv="us.img.e-planning.net" data-sv="ads.us.e-planning.net" data-ci="1dc9a" data-usedivname="true"></script>

<script>
(function (ci) {
  var x, o = window.document, s = (o.location.protocol=="https:"), h = o.createElement("script"), d = "e-planning.net", i = (s?"us":"aklc")+".img."+d;
  var a = {"data-isv": i, "data-sv":"ads.us."+d, "data-ci":ci, id:"hbepl", async:"async", src:"http"+(s?"s":"")+"://"+i+"/layers/hbdfp.js"};
  for (x in a) 
    h.setAttribute(x, a[x]);
  o.head.appendChild(h);
})("1dc9a");
</script>
-->

<script type='text/javascript'>
zonaTO = 'Portada';
var ct_prog = [""];
var ct_seccion = ["home"];
         
var googletag = googletag || {};
googletag.cmd = googletag.cmd || [];
(function() {
	var gads = document.createElement('script');
	gads.async = true;
	gads.type = 'text/javascript';
	var useSSL = 'https:' == document.location.protocol;
	gads.src = (useSSL ? 'https:' : 'http:') + 
	'//www.googletagservices.com/tag/js/gpt.js';
	var node = document.getElementsByTagName('script')[0];
	node.parentNode.insertBefore(gads, node);
})();
</script>
<script type='text/javascript'>
portada=0;
googletag.cmd.push(function() {
   /**
var mapBanner = googletag.sizeMapping().
		addSize([320, 400], [320, 50]).
        addSize([320, 568], [320, 50]).
        addSize([980, 690], [728, 90]).
		addSize([1024, 768], [970,90]).
		addSize([1024, 768], [728,90]).
		build();
**/

if (deviceDetect() != 'mobile' ){
        googletag.defineSlot('/148773018/Canal12_ROS', [[728, 90], [960, 90]], 'div-gpt-ad-topbanner').
        addService(googletag.companionAds()).addService(googletag.pubads());
        googletag.defineSlot('/148773018/Canal12_ROS', [[728, 90], [960, 90]], 'div-gpt-ad-midbanner').
        addService(googletag.companionAds()).addService(googletag.pubads());
        googletag.defineSlot('/148773018/Canal12_ROS', [[300, 250]], 'div-gpt-ad-boton').
        addService(googletag.companionAds()).addService(googletag.pubads());
        googletag.defineOutOfPageSlot('/148773018/Canal12_ROS', 'div-gpt-ad-oop').addService(googletag.pubads()).setTargeting("pos", "inter");
    }else{
        googletag.defineSlot('/148773018/Canal12_ROS', [[320, 50]], 'div-gpt-ad-topbanner').
        addService(googletag.companionAds()).addService(googletag.pubads());
        googletag.defineSlot('/148773018/Canal12_ROS', [[320, 50]], 'div-gpt-ad-midbanner').
        addService(googletag.companionAds()).addService(googletag.pubads());
        googletag.defineSlot('/148773018/Canal12_ROS', [[300, 250]], 'div-gpt-ad-boton').
        addService(googletag.companionAds()).addService(googletag.pubads());
    }

	googletag.pubads().setTargeting("ct_seccion", ct_seccion);
	googletag.pubads().enableSingleRequest();
	googletag.pubads().collapseEmptyDivs(true);
	googletag.enableServices();
});
</script>
</head>
<body data-ga="Home" data-ga-seccion="Principal" data-ga-id="home">
<div id="fb-root"></div>
<script type="text/javascript">
    rutacc = '';
</script>
<script>
(function(d, s, id) {
  var js, fjs = d.getElementsByTagName(s)[0];
  if (d.getElementById(id)) return;
  js = d.createElement(s); js.id = id;
  js.src = "//connect.facebook.net/es_LA/sdk.js#xfbml=1&appId=782051041914141&version=v2.3";
  fjs.parentNode.insertBefore(js, fjs);
}(document, 'script', 'facebook-jssdk'));
</script>
<script>
  (function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
  (i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
  m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
  })(window,document,'script','//www.google-analytics.com/analytics.js','ga');

  ga('create', 'UA-5745109-2', 'auto');
  
  if (typeof autor_nodo != 'undefined'){
      ga('set', 'dimension1', autor_nodo);
  }
  if (typeof origen_nodo != 'undefined'){
      if (autor_nodo == "ned") origen_nodo = "NED: " + origen_nodo;
      ga('set', 'dimension2', origen_nodo);
  }

  if (typeof tagList != 'undefined' && tagList.length > 0) {
      for (i = 0; i < tagList.length; i++) {
          ga('set', 'dimension3', tagList[i]);
      }
  }

  ga('send', 'pageview');
</script>
<script src="http://cdn.canal12.com.sv/sites/common/js/tracking.js"></script>
<script async src="https://cdn.onthe.io/io.js/YcJ0UhfdeXpu"></script>
<header id="headerTop">
  <div id="banner">
    <div id="zonaPushdown">
      <div id="pushdown"></div>
    </div>
  </div>
</header>
<nav id="menumobile">
  <div class="icomenu" data-toggle="modal" data-target="#modalMenu"></div>
  <a href="/" class="icologo"></a> <a href="/contactenos" class="contact"></a>
  <div class="search"></div>
  <a href="/envivo" id="envivo"> <span class="cab">
  <div class="ico"></div>
  <div class="desc">en vivo</div>
  </span> </a>
  <div id="modalmobile">
    <div class="cerrar">[x]cerrar</div>
    <div id="menuint">
      <ul>
        <li><a href="/noticias/actualidad-1">Actualidad</a></li>
        <li><a href="/noticias/deportes-3">Deportes</a></li>
        <li><a href="/noticias/espectaculos-2">Espectáculos</a></li>
        <li><a href="/noticias">Noticias</a></li>
        <li><a href="/programas">Programas</a></li>
        <li><a href="/novelas">Novelas</a></li>
        <li><a href="/envivo">En Vivo</a></li>
      </ul>
    </div>
  </div>
</nav>
<div id="searchmobile">
  <input type="text" class="buscador" placeholder="buscar...">
  <div class="ico"></div>
</div>
<section id="slideshow" class="homeslideshow">
  <nav id="menumain">
  <ul>
    <li class="dditem" id="itm_menu">
      <div class="ico"></div>
      <span>MENU</span>
      <ul class="ddmenu">
        <li><a href="/noticias/actualidad-1">Actualidad</a></li>
        <li><a href="/noticias/deportes-3">Deportes</a></li>
        <li><a href="/noticias/espectaculos-2">Espectáculos</a></li>
        <li><a href="/noticias">Noticias</a></li>
        <li><a href="/programas">Programas</a></li>
        <li><a href="/novelas">Novelas</a></li>
        <li><a href="/envivo">En Vivo</a></li>
      </ul>
    </li>
    <li class="logoMain"><a href="/"></a></li>
    <li class="itmseccion"><a href="/noticias">NOTICIAS</a></li>
    <li class="itmseccion"><a  href="/noticias/actualidad-1">ACTUALIDAD</a></li>
    <li class="itmseccion"><a  href="/noticias/deportes-3">DEPORTES</a></li>
    <li class="itmseccion"><a  href="/noticias/espectaculos-2">ESPECTÁCULOS</a></li>
    <li class="dditem" id="itm_programas"><a href="/programas">PROGRAMAS</a>
      <div class="icodown"></div>
      <ul class="ddmenu">
        <li><a href="/programa/cinema-12">Cinema 12</a></li>
        <li><a href="/programa/hola-el-salvador">Hola El Salvador</a></li>
        <li><a href="/programa/noticiero-hechos-estelar">Noticiero Hechos Estelar</a></li>
        <li><a href="/programa/pizarron-deportivo">Pizarrón Deportivo</a></li>
        <li><a href="/programa/pop-12">Pop 12</a></li>
        <li><a href="/programas">Más Programas</a></li>
      </ul>
    </li>
    <li class="dditem" id="itm_novelas"><a href="/novelas">NOVELAS</a>
      <div class="icodown"></div>
      <ul class="ddmenu">
        <li><a href="/programa/a-cada-quien-su-santo">A Cada Quien Su Santo</a></li>
        <li><a href="/programa/cambio-de-vida">Cambio de Vida</a></li>
        <li><a href="/novelas">Más Novelas</a></li>
      </ul>
    </li>
    <li class="dditem" id="itm_series"><a href="/series">SERIES</a>
      <div class="icodown"></div>
      <ul class="ddmenu">
        <li><a href="/series">Más Series</a></li>
      </ul>
    </li>
    <li class="dditem" id="itm_paises"><a style="padding-right: 2px; color:rgba(255,255,255,0.5);">PAIS</a>
      <div class="escudo_pais el_salvador"></div>
      <div class="icodown paises"></div>
      <ul class="ddmenu paises">
        <li class="paises"><a href="http://www.elnueve.com.ar" class="paises" target="_blank">
          <div class="izquierda">Argentina</div>
          <div class="derecha">
            <div class="escudo_pais argentina"></div>
          </div>
          </a></li>
          <li class="paises"><a href="http://www.redbolivision.tv.bo" class="paises" target="_blank">
          <div class="izquierda">Bolivia</div>
          <div class="derecha">
            <div class="escudo_pais bolivia"></div>
          </div>
          </a></li>
        <li class="paises"><a href="http://www.repretel.com" class="paises" target="_blank">
          <div class="izquierda">Costa Rica</div>
          <div class="derecha">
            <div class="escudo_pais costa_rica"></div>
          </div>
          </a></li>
        <li class="paises smi">
          <div class="sub-menu1">
            <div class="izquierda">Ecuador</div>
            <div class="derecha">
              <div class="escudo_pais ecuador"></div>
            </div>
            <ul class="sub-menu2">
              <li class="paises"> <a href="http://www.rts.com.ec" class="paises" target="_blank">
                <div class="izquierda">RTS</div>
                <div class="derecha"> <img src="http://cdn.rts.com.ec/sites/common/img/logo_rts.png" height="20" /> </div>
                </a> </li>
              <li class="paises"> <a href="http://www.tvc.com.ec" class="paises" target="_blank">
                <div class="izquierda">TVC</div>
                <div class="derecha"> <img src="http://cdn.tvc.com.ec/sites/common/img/logo_televicentro.png" height="20" /> </div>
                </a> </li>
            </ul>
          </div>
        </li>
        <li class="paises"><a href="http://www.chapintv.com" class="paises" target="_blank">
          <div class="izquierda">Guatemala</div>
          <div class="derecha">
            <div class="escudo_pais guatemala"></div>
          </div>
          </a></li>
        <li class="paises"><a href="http://www.vtv.com.hn" class="paises" target="_blank">
          <div class="izquierda">Honduras</div>
          <div class="derecha">
            <div class="escudo_pais honduras"></div>
          </div>
          </a></li>
        <li class="paises"><a href="http://www.canal10.com.ni" class="paises" target="_blank">
          <div class="izquierda">Nicaragua</div>
          <div class="derecha">
            <div class="escudo_pais nicaragua"></div>
          </div>
          </a></li>
        <li class="paises"><a href="http://www.snt.com.py" class="paises" target="_blank">
          <div class="izquierda">Paraguay</div>
          <div class="derecha">
            <div class="escudo_pais paraguay"></div>
          </div>
          </a></li>
        <li class="paises smi">
          <div class="sub-menu1">
            <div class="izquierda">Perú</div>
            <div class="derecha">
              <div class="escudo_pais peru"></div>
            </div>
            <ul class="sub-menu2">
              <li class="paises"> <a href="http://www.atv.pe" class="paises" target="_blank">
                <div class="izquierda">ATV</div>
                <div class="derecha"> <img src="http://cdn.atv.pe/sites/atv.pe/common/img/logo_atvpe.png" height="20" /> </div>
                </a> </li>
            </ul>
          </div>
        </li>
        <li class="paises"><a href="http://www.antena7.com.do" class="paises" target="_blank">
          <div class="izquierda">Rep. Dom.</div>
          <div class="derecha">
            <div class="escudo_pais republica_dominicana"></div>
          </div>
          </a></li>
      </ul>
    </li>
    <li style="padding-top: 12px; position: relative; padding-left: 2px">
      <input type="text" id="buscadorTop" class="buscador"  />
      <div class="iconobusc"></div>
    </li>
    <li class="dditem" style="padding-top: 11px" id="itm_canales"> <a id="envivo" href="/envivo"> <span class="cab">
      <div class="ico"></div>
      <div class="desc">en vivo</div>
      </span> </a>
    </li>
  </ul>
</nav>
  
<div id="carousel-slide" class="carousel slide" data-ride="carousel"> 
  <!-- Indicators -->
  <ol class="carousel-indicators">
        <li data-target="#carousel-slide" data-slide-to="0" class="active"></li>
        <li data-target="#carousel-slide" data-slide-to="1" ></li>
      </ol>
  
  <!-- Wrapper for slides -->
  <div class="carousel-inner home" id="lista">
        <div class="item active" style="background-image:url(http://cdn.canal12.com.sv/files/2018/03/20/banner-01_.jpg);">
    <a href="http://www.canal12.com.sv/actualidad/blind-2-chat-51777" style="width:100%; height:100%; position:absolute;">
      <div class="layer anuncio" style="width: 100%;"></div>
      <div class="desc"> 
                        <h1>Blind 2 Chat</h1>
        <h2></h2>
        <div class="tags" style="display:none;">
                            </div>
      </div>
        </a>
    </div>
        <div class="item " style="background-image:url(http://cdn.canal12.com.sv/files/2017/08/22/web-Rosa-Negra-Banner-Miralo.jpg);">
    <a href="http://www.canal12.com.sv/actualidad/rosa-negra-36303" style="width:100%; height:100%; position:absolute;">
      <div class="layer " style="width: 100%;"></div>
      <div class="desc"> 
                        <h1>Rosa Negra</h1>
        <h2>Lunes A Viernes (6:00 pm - 7:00 pm) por Canal 12</h2>
        <div class="tags" style="display:none;">
                            </div>
      </div>
        </a>
    </div>
      </div>
  
  <!-- Controls --> 
  <a class="left carousel-control" href="#carousel-slide" role="button" data-slide="prev"> <span class="botnav prev"></span> </a> <a class="right carousel-control" href="#carousel-slide" role="button" data-slide="next"> <span class="botnav next"></span> </a> </div>
  <div class="pie home">
    <div class="cont"> </div>
  </div>
  <div class="shadowpie"></div>
</section>
<section id="main" class="contenedor" >
  <div id="bloqueredes">
    <ul>
      <li>
        <div class="fb-like" data-href="http://www.facebook.com/CanalDoceSV" data-layout="button_count" data-action="like" data-show-faces="false" data-share="true"></div>
      </li>
      <li><a class="twitter-follow-button" href="http://www.twitter.com/Canal_12" data-show-count="true" data-lang="es"> Sigue @Canal_12 </a> 
        <script type="text/javascript">
window.twttr = (function (d, s, id) {
  var t, js, fjs = d.getElementsByTagName(s)[0];
  if (d.getElementById(id)) return;
  js = d.createElement(s); js.id = id;
  js.src= "https://platform.twitter.com/widgets.js";
  fjs.parentNode.insertBefore(js, fjs);
  return window.twttr || (t = { _e: [], ready: function (f) { t._e.push(f) } });
}(document, "script", "twitter-wjs"));
</script></li>
      <li><!-- Place this tag in your head or just before your close body tag. --> 
        <script src="https://apis.google.com/js/platform.js" async defer>
  {lang: 'es-419'}
</script> 
        
        <!-- Place this tag where you want the widget to render. -->
        <div class="g-follow" data-annotation="bubble" data-height="20" data-href="http://plus.google.com/100912321241699444897" data-rel="publisher"></div>
      </li>
    </ul>
    <div class="texto">Síguenos en nuestras redes</div>
  </div>
  <section id="programacion">
    <div class="cab">PROGRAMACIÓN <span>Canal 12</span></div>
      <!-- Indicators -->
 
  <div class="" id="listaini">
        <a href="http://www.canal12.com.sv/envivo" class="item itemrel active"><img data-original="http://cdn.canal12.com.sv/files/2017/04/26/320x150_rosa-negras-mantenimiento.jpg" class="lazy" alt="Rosa Negra" title="Rosa Negra" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/04/26/320x150_rosa-negras-mantenimiento.jpg" alt="Rosa Negra" title="Rosa Negra" /></noscript>
    <div class="info"> <span class="ahora">ahora</span> <b> 18:00 h</b><br>
      <span class="ht">Rosa Negra</span><br>
      <span class="lv">Lunes a Viernes</span> </div>
    </a>
        <a href="#" class="item itemrel sec"><img data-original="http://cdn.canal12.com.sv/files/2018/01/15/320x150_feriha_0.jpg" class="lazy" alt="El Secreto de Feriha" title="El Secreto de Feriha" /><noscript><img src="http://cdn.canal12.com.sv/files/2018/01/15/320x150_feriha_0.jpg" alt="El Secreto de Feriha" title="El Secreto de Feriha" /></noscript>
    <div class="info"> <span class="">a continuación</span> <b> 19:00 h</b><br>
      <span class="ht">El Secreto de Feriha</span><br>
      <span class="lv">Lunes a Viernes</span> </div>
    </a>
        <a href="#" class="item itemrel sec"><img data-original="http://cdn.canal12.com.sv/files/2017/03/08/hechos-estelar_0.jpg" class="lazy" alt="Noticiero Hechos Estelar" title="Noticiero Hechos Estelar" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/03/08/hechos-estelar_0.jpg" alt="Noticiero Hechos Estelar" title="Noticiero Hechos Estelar" /></noscript>
    <div class="info"> <span class="">después</span> <b> 20:00 hrs</b><br>
      <span class="ht">Noticiero Hechos Estelar</span><br>
      <span class="lv">Lunes a Viernes</span> </div>
    </a>
      </div>
  </section>
  <section id="listapastillas" class="nomask">
    <div class="cab">
      <div style="float:left">VIDEOS</div>
      <div style="float:right"><script src="https://apis.google.com/js/platform.js"></script>
        <div class="g-ytsubscribe" data-channel="canal12sv" data-layout="default" data-count="undefined"></div>
      </div>
    </div>
    <div class="lista">
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/mostramos-principales-novedades-cinematograficas-51836">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_25.612Z_image.jpg" class="img_def lazy" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_25.612Z_image.jpg" class="img_def" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_25.612Z_image.jpg" class="img_small lazy" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_25.612Z_image.jpg" class="img_small" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_25.612Z_image.jpg" class="img_tiny lazy" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_25.612Z_image.jpg" class="img_tiny" alt="Le mostramos las principales novedades cinematográficas" title="Le mostramos las principales novedades cinematográficas"></noscript>
          <div class="titulo">Le mostramos las principales novedades cinematográficas</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/mostramos-principales-novedades-cinematograficas-51836"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/mostramos-principales-novedades-cinematograficas-51836" sharetext="Le mostramos las principales novedades cinematográficas via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/mostramos-principales-novedades-cinematograficas-51836"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/delicias-culinarias-preparamos-sabrosas-pechugas-rellenas-vegetales-51835">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_24.950Z_image.jpg" class="img_def lazy" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_24.950Z_image.jpg" class="img_def" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_24.950Z_image.jpg" class="img_small lazy" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_24.950Z_image.jpg" class="img_small" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_24.950Z_image.jpg" class="img_tiny lazy" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_24.950Z_image.jpg" class="img_tiny" alt="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''" title="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''"></noscript>
          <div class="titulo">Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales''</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/delicias-culinarias-preparamos-sabrosas-pechugas-rellenas-vegetales-51835"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/delicias-culinarias-preparamos-sabrosas-pechugas-rellenas-vegetales-51835" sharetext="Delicias culinarias: Preparamos unas sabrosas ''pechugas rellenas de vegetales'' via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/delicias-culinarias-preparamos-sabrosas-pechugas-rellenas-vegetales-51835"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/increible-parezca-piscina-puede-desaparecer-cosa-minutos-51834">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_24.514Z_image.jpg" class="img_def lazy" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_24.514Z_image.jpg" class="img_def" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_24.514Z_image.jpg" class="img_small lazy" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_24.514Z_image.jpg" class="img_small" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_24.514Z_image.jpg" class="img_tiny lazy" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_24.514Z_image.jpg" class="img_tiny" alt="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos" title="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos"></noscript>
          <div class="titulo">Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/increible-parezca-piscina-puede-desaparecer-cosa-minutos-51834"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/increible-parezca-piscina-puede-desaparecer-cosa-minutos-51834" sharetext="Por Increíble que parezca: Piscina puede desaparecer en cosa de minutos via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/increible-parezca-piscina-puede-desaparecer-cosa-minutos-51834"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/rene-rivas-habla-sobre-exito-youtube-51833">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_23.305Z_image.jpg" class="img_def lazy" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_23.305Z_image.jpg" class="img_def" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_23.305Z_image.jpg" class="img_small lazy" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_23.305Z_image.jpg" class="img_small" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_23.305Z_image.jpg" class="img_tiny lazy" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_23.305Z_image.jpg" class="img_tiny" alt="René Rivas nos habla sobre su éxito en YouTube" title="René Rivas nos habla sobre su éxito en YouTube"></noscript>
          <div class="titulo">René Rivas nos habla sobre su éxito en YouTube</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/rene-rivas-habla-sobre-exito-youtube-51833"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/rene-rivas-habla-sobre-exito-youtube-51833" sharetext="René Rivas nos habla sobre su éxito en YouTube via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/rene-rivas-habla-sobre-exito-youtube-51833"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/cinco-cosas-debe-hacer-padre-hijos-51832">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_22.416Z_image.jpg" class="img_def lazy" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_22.416Z_image.jpg" class="img_def" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_22.416Z_image.jpg" class="img_small lazy" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_22.416Z_image.jpg" class="img_small" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_22.416Z_image.jpg" class="img_tiny lazy" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_22.416Z_image.jpg" class="img_tiny" alt="Estas son las cinco cosas que debe hacer un padre por sus hijos" title="Estas son las cinco cosas que debe hacer un padre por sus hijos"></noscript>
          <div class="titulo">Estas son las cinco cosas que debe hacer un padre por sus hijos</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/cinco-cosas-debe-hacer-padre-hijos-51832"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/cinco-cosas-debe-hacer-padre-hijos-51832" sharetext="Estas son las cinco cosas que debe hacer un padre por sus hijos via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/cinco-cosas-debe-hacer-padre-hijos-51832"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/conmemora-dia-mundial-sindrome-down-51830">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_21.196Z_image.jpg" class="img_def lazy" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_21.196Z_image.jpg" class="img_def" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_21.196Z_image.jpg" class="img_small lazy" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_21.196Z_image.jpg" class="img_small" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_21.196Z_image.jpg" class="img_tiny lazy" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_21.196Z_image.jpg" class="img_tiny" alt="Hoy se conmemora el ''Día Mundial del Síndrome de Down''" title="Hoy se conmemora el ''Día Mundial del Síndrome de Down''"></noscript>
          <div class="titulo">Hoy se conmemora el ''Día Mundial del Síndrome de Down''</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/conmemora-dia-mundial-sindrome-down-51830"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/conmemora-dia-mundial-sindrome-down-51830" sharetext="Hoy se conmemora el ''Día Mundial del Síndrome de Down'' via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/conmemora-dia-mundial-sindrome-down-51830"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/revisamos-publicaciones-importantes-redes-sociales-51827">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_19.962Z_image.jpg" class="img_def lazy" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_19.962Z_image.jpg" class="img_def" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_19.962Z_image.jpg" class="img_small lazy" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_19.962Z_image.jpg" class="img_small" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_19.962Z_image.jpg" class="img_tiny lazy" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_19.962Z_image.jpg" class="img_tiny" alt="Revisamos las publicaciones más importantes en las redes sociales" title="Revisamos las publicaciones más importantes en las redes sociales"></noscript>
          <div class="titulo">Revisamos las publicaciones más importantes en las redes sociales</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/revisamos-publicaciones-importantes-redes-sociales-51827"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/revisamos-publicaciones-importantes-redes-sociales-51827" sharetext="Revisamos las publicaciones más importantes en las redes sociales via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/revisamos-publicaciones-importantes-redes-sociales-51827"></div>
            </div>
          </div>
        </div>
  
     <div class="item "> <a href="http://www.canal12.com.sv/actualidad/negocios-hechos-empresas-buscan-personal-domine-diversos-idiomas-51825">
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_16.736Z_image.jpg" class="img_def lazy" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/2018-03-21T12_20_16.736Z_image.jpg" class="img_def" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_16.736Z_image.jpg" class="img_small lazy" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/316x202_2018-03-21T12_20_16.736Z_image.jpg" class="img_small" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas"></noscript>
     <img data-original="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_16.736Z_image.jpg" class="img_tiny lazy" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas">
     <noscript><img src="http://cdn.canal12.com.sv/files/2018/03/21/175x112_2018-03-21T12_20_16.736Z_image.jpg" class="img_tiny" alt="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas" title="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas"></noscript>
          <div class="titulo">Negocios Hechos: Empresas buscan a personal que domine diversos idiomas</div>
          </a>
          <div class="redes"><span>Compartir en:</span>
            <div class="list">
              <div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/actualidad/negocios-hechos-empresas-buscan-personal-domine-diversos-idiomas-51825"></div>
              <div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/actualidad/negocios-hechos-empresas-buscan-personal-domine-diversos-idiomas-51825" sharetext="Negocios Hechos: Empresas buscan a personal que domine diversos idiomas via @#"></div>
              <div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/actualidad/negocios-hechos-empresas-buscan-personal-domine-diversos-idiomas-51825"></div>
            </div>
          </div>
        </div>
    
</div>
  </section>
  <section id="listaprogramas">
    <div class="cab">PROGRAMAS</div>
    <div class="mask">
      <div class="lista">
    <a href="http://www.canal12.com.sv/programa/cinema-12"> <img data-original="http://cdn.canal12.com.sv/files/2017/08/09/188x265_cinema12_0.jpg" class="lazy" alt="Cinema 12" title="Cinema 12" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/08/09/188x265_cinema12_0.jpg" alt="Cinema 12" title="Cinema 12" /></noscript>
  <div class="titulo">Cinema 12</div>
  </a>
    <a href="http://www.canal12.com.sv/programa/pizarron-deportivo"> <img data-original="http://cdn.canal12.com.sv/files/2017/11/01/188x265_plantilla_pdnoche.jpg" class="lazy" alt="Pizarrón Deportivo" title="Pizarrón Deportivo" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/11/01/188x265_plantilla_pdnoche.jpg" alt="Pizarrón Deportivo" title="Pizarrón Deportivo" /></noscript>
  <div class="titulo">Pizarrón Deportivo</div>
  </a>
    <a href="http://www.canal12.com.sv/programa/pop-12"> <img data-original="http://cdn.canal12.com.sv/files/2017/03/10/188x265_pop-12.jpg" class="lazy" alt="Pop 12" title="Pop 12" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/03/10/188x265_pop-12.jpg" alt="Pop 12" title="Pop 12" /></noscript>
  <div class="titulo">Pop 12</div>
  </a>
  </div>
    </div>
  </section>
  <hr>
  <section id="listanovelas">
    <div class="cab">NOVELAS</div>
    <div class="mask">
      <div class="lista">
    <a href="http://www.canal12.com.sv/programa/esperanza-el-destino-del-amor"> <img data-original="http://cdn.canal12.com.sv/files/2018/01/18/188x265_esperanza_0.jpg" class="lazy" alt="Esperanza, el destino del amor" title="Esperanza, el destino del amor" /><noscript><img src="http://cdn.canal12.com.sv/files/2018/01/18/188x265_esperanza_0.jpg" alt="Esperanza, el destino del amor" title="Esperanza, el destino del amor" /></noscript>
  <div class="titulo">Esperanza, el destino del amor</div>
  </a>
    <a href="http://www.canal12.com.sv/programa/rosa-negra"> <img data-original="http://cdn.canal12.com.sv/files/2017/04/26/188x265_rosa-negra_0.jpg" class="lazy" alt="Rosa Negra" title="Rosa Negra" /><noscript><img src="http://cdn.canal12.com.sv/files/2017/04/26/188x265_rosa-negra_0.jpg" alt="Rosa Negra" title="Rosa Negra" /></noscript>
  <div class="titulo">Rosa Negra</div>
  </a>
    <a href="#"> <img data-original="" class="lazy" alt="El Secreto de Feriha" title="El Secreto de Feriha" /><noscript><img src="" alt="El Secreto de Feriha" title="El Secreto de Feriha" /></noscript>
  <div class="titulo">El Secreto de Feriha</div>
  </a>
    <a href="http://www.canal12.com.sv/programa/sila"> <img data-original="http://cdn.canal12.com.sv/files/2018/01/15/188x265_sila_0.jpg" class="lazy" alt="Sila" title="Sila" /><noscript><img src="http://cdn.canal12.com.sv/files/2018/01/15/188x265_sila_0.jpg" alt="Sila" title="Sila" /></noscript>
  <div class="titulo">Sila</div>
  </a>
    <a href="http://www.canal12.com.sv/programa/a-cada-quien-su-santo"> <img data-original="http://cdn.canal12.com.sv/files/2015/12/08/a_cada_quien_su_santo_.jpg" class="lazy" alt="A Cada Quien su Santo" title="A Cada Quien su Santo" /><noscript><img src="http://cdn.canal12.com.sv/files/2015/12/08/a_cada_quien_su_santo_.jpg" alt="A Cada Quien su Santo" title="A Cada Quien su Santo" /></noscript>
  <div class="titulo">A Cada Quien su Santo</div>
  </a>
  </div>
    </div>
  </section>
  <section id="bannermedio">
    <!-- /midbanner/Canal_9 -->
<div id='div-gpt-ad-midbanner' class="adunit_standard">
<script type='text/javascript'>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-midbanner'); });
</script>
</div>  </section>
  <section id="lafrase">
    <div class="cab"><span>LA FRASE</span>
      <div class="ico"></div>
    </div>
    <svg width="22" height="54" style="float: left" >
    <polygon points="0,0,22,27,0,54" style="fill:black;stroke:black;stroke-width:0" />
    </svg>
    <div class="cont">
	<span>"No teníamos conocimiento que Gustavito estuviera enfermo"<a href="http://www.canal12.com.sv/actualidad/secretaria-cultura-entrega-declaracion-por-muerte-gustavito-33692" class="botonenlace botlink" style="margin-left:5px">ir a la noticia</a></span>
</div>  </section>
  <table class="bloquenotas" id="bloqueNotas1">
	<tr>
		<td id="columna_1"><article class="item" id="article_1_1">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/el-momento-en-que-una-mujer-da-a-luz-mientras-se-bana-en-el-mar-51474">
					<h2>El momento en que una mujer da a luz mientras se baña en el mar</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/el-momento-en-que-una-mujer-da-a-luz-mientras-se-bana-en-el-mar-51474"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/el-momento-en-que-una-mujer-da-a-luz-mientras-se-bana-en-el-mar-51474" sharetext="El momento en que una mujer da a luz mientras se baña en el mar #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/el-momento-en-que-una-mujer-da-a-luz-mientras-se-bana-en-el-mar-51474"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/el-momento-en-que-una-mujer-da-a-luz-mientras-se-bana-en-el-mar-51474">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa80c997411f51a58ef3ef6.jpg" class="img_def lazy" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa80c997411f51a58ef3ef6.jpg" class="img_def" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa80c997411f51a58ef3ef6.jpg" class="img_small lazy" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa80c997411f51a58ef3ef6.jpg" class="img_small" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa80c997411f51a58ef3ef6.jpg" class="img_tiny lazy" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa80c997411f51a58ef3ef6.jpg" class="img_tiny" alt="El momento en que una mujer da a luz mientras se baña en el mar" title="El momento en que una mujer da a luz mientras se baña en el mar"></noscript>
					</div>
    				<h3>El insólito hecho fue captado en el balneario de Dahab en el Mar Rojo en Egipto.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_3">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/asistio-a-300-conciertos-de-luis-miguel-y-recibio-un-premio-inesperado-de-parte-del-artista-51471">
					<h2>Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/asistio-a-300-conciertos-de-luis-miguel-y-recibio-un-premio-inesperado-de-parte-del-artista-51471"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/asistio-a-300-conciertos-de-luis-miguel-y-recibio-un-premio-inesperado-de-parte-del-artista-51471" sharetext="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/asistio-a-300-conciertos-de-luis-miguel-y-recibio-un-premio-inesperado-de-parte-del-artista-51471"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/asistio-a-300-conciertos-de-luis-miguel-y-recibio-un-premio-inesperado-de-parte-del-artista-51471">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa7ea4b7411f51a58ef391e.jpg" class="img_def lazy" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa7ea4b7411f51a58ef391e.jpg" class="img_def" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa7ea4b7411f51a58ef391e.jpg" class="img_small lazy" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa7ea4b7411f51a58ef391e.jpg" class="img_small" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa7ea4b7411f51a58ef391e.jpg" class="img_tiny lazy" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa7ea4b7411f51a58ef391e.jpg" class="img_tiny" alt="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista" title="Asistió a 300 conciertos de Luis Miguel y recibió un premio inesperado de parte del artista"></noscript>
					</div>
    				<h3>"El Sol de México" advirtió la presencia de la mujer en el público, en pleno show, y se acercó a ella.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_6">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/ken-humano-muestra-las-costillas-que-le-quitaron-y-sus-seguidores-exigen-que-elimine-la-foto-51393">
					<h2>"Ken Humano" muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/ken-humano-muestra-las-costillas-que-le-quitaron-y-sus-seguidores-exigen-que-elimine-la-foto-51393"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/ken-humano-muestra-las-costillas-que-le-quitaron-y-sus-seguidores-exigen-que-elimine-la-foto-51393" sharetext=""Ken Humano" muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/ken-humano-muestra-las-costillas-que-le-quitaron-y-sus-seguidores-exigen-que-elimine-la-foto-51393"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/ken-humano-muestra-las-costillas-que-le-quitaron-y-sus-seguidores-exigen-que-elimine-la-foto-51393">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa680fe7411f50fa7c6fa5e.jpg" class="img_def lazy" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa680fe7411f50fa7c6fa5e.jpg" class="img_def" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa680fe7411f50fa7c6fa5e.jpg" class="img_small lazy" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa680fe7411f50fa7c6fa5e.jpg" class="img_small" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa680fe7411f50fa7c6fa5e.jpg" class="img_tiny lazy" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa680fe7411f50fa7c6fa5e.jpg" class="img_tiny" alt="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto" title="Ken Humano muestra las costillas que le quitaron y sus seguidores exigen que elimine la foto"></noscript>
					</div>
    				<h3>Cientos de críticas recibió, luego de publicar la polémica imagen que perturbó a sus seguidores.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_9">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/cuanto-te-costaria-clonar-a-tu-mascota-50963">
					<h2>¿Cuánto te costaría clonar a tu mascota?</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/cuanto-te-costaria-clonar-a-tu-mascota-50963"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/cuanto-te-costaria-clonar-a-tu-mascota-50963" sharetext="¿Cuánto te costaría clonar a tu mascota? #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/cuanto-te-costaria-clonar-a-tu-mascota-50963"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/cuanto-te-costaria-clonar-a-tu-mascota-50963">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5a97fb907411f553d721847e.jpg" class="img_def lazy" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?">
						<noscript><img src="http://cdn.canal12.com.sv/files/5a97fb907411f553d721847e.jpg" class="img_def" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5a97fb907411f553d721847e.jpg" class="img_small lazy" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5a97fb907411f553d721847e.jpg" class="img_small" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5a97fb907411f553d721847e.jpg" class="img_tiny lazy" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5a97fb907411f553d721847e.jpg" class="img_tiny" alt="¿Cuánto te costaría clonar a tu mascota?" title="¿Cuánto te costaría clonar a tu mascota?"></noscript>
					</div>
    				<h3>En Estados Unidos hay una empresa que se dedica a prestar este servicio, el que por supuesto no es nada barato.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article></td>
		<td id="columna_2"><article class="item" id="article_1_2">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/el-perro-con-rostro-humano-que-desata-la-locura-de-los-usuarios-en-la-web-51462">
					<h2>El perro con "rostro humano" que desata la locura de los usuarios en la web</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/el-perro-con-rostro-humano-que-desata-la-locura-de-los-usuarios-en-la-web-51462"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/el-perro-con-rostro-humano-que-desata-la-locura-de-los-usuarios-en-la-web-51462" sharetext="El perro con "rostro humano" que desata la locura de los usuarios en la web #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/el-perro-con-rostro-humano-que-desata-la-locura-de-los-usuarios-en-la-web-51462"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/el-perro-con-rostro-humano-que-desata-la-locura-de-los-usuarios-en-la-web-51462">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa7eb1e7411f51a58ef3983.jpg" class="img_def lazy" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa7eb1e7411f51a58ef3983.jpg" class="img_def" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa7eb1e7411f51a58ef3983.jpg" class="img_small lazy" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa7eb1e7411f51a58ef3983.jpg" class="img_small" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa7eb1e7411f51a58ef3983.jpg" class="img_tiny lazy" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa7eb1e7411f51a58ef3983.jpg" class="img_tiny" alt="El perro con rostro humano que desata la locura de los usuarios en la web" title="El perro con rostro humano que desata la locura de los usuarios en la web"></noscript>
					</div>
    				<h3>La inquietante apariencia del animal hizo que su foto se viralizara en las redes sociales.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_4">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/llego-a-su-fin-la-extrana-batalla-legal-por-el-cadaver-de-charles-manson -51468">
					<h2>Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson </h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/llego-a-su-fin-la-extrana-batalla-legal-por-el-cadaver-de-charles-manson -51468"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/llego-a-su-fin-la-extrana-batalla-legal-por-el-cadaver-de-charles-manson -51468" sharetext="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson  #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/llego-a-su-fin-la-extrana-batalla-legal-por-el-cadaver-de-charles-manson -51468"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/llego-a-su-fin-la-extrana-batalla-legal-por-el-cadaver-de-charles-manson -51468">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa7fdd97411f51a58ef3ca4.jpg" class="img_def lazy" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson ">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa7fdd97411f51a58ef3ca4.jpg" class="img_def" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson "></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa7fdd97411f51a58ef3ca4.jpg" class="img_small lazy" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson ">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa7fdd97411f51a58ef3ca4.jpg" class="img_small" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson "></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa7fdd97411f51a58ef3ca4.jpg" class="img_tiny lazy" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson ">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa7fdd97411f51a58ef3ca4.jpg" class="img_tiny" alt="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson " title="Llegó a su fin la extraña batalla legal por el cadáver de Charles Manson "></noscript>
					</div>
    				<h3>La Corte Superior de Kern confirmó que el cuerpo será entregado a un nieto del psicópata.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_7">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/fue-a-una-fiesta-vio-a-su-novia-besandose-con-otro-y-su-inesperada-reaccion-se-hizo-viral-51407">
					<h2>Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/fue-a-una-fiesta-vio-a-su-novia-besandose-con-otro-y-su-inesperada-reaccion-se-hizo-viral-51407"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/fue-a-una-fiesta-vio-a-su-novia-besandose-con-otro-y-su-inesperada-reaccion-se-hizo-viral-51407" sharetext="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/fue-a-una-fiesta-vio-a-su-novia-besandose-con-otro-y-su-inesperada-reaccion-se-hizo-viral-51407"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/fue-a-una-fiesta-vio-a-su-novia-besandose-con-otro-y-su-inesperada-reaccion-se-hizo-viral-51407">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa6a9f47411f50fa7c7036f.jpg" class="img_def lazy" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa6a9f47411f50fa7c7036f.jpg" class="img_def" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa6a9f47411f50fa7c7036f.jpg" class="img_small lazy" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa6a9f47411f50fa7c7036f.jpg" class="img_small" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa6a9f47411f50fa7c7036f.jpg" class="img_tiny lazy" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa6a9f47411f50fa7c7036f.jpg" class="img_tiny" alt="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral" title="Fue a una fiesta, vio a su novia besándose con otro y su inesperada reacción se hizo viral"></noscript>
					</div>
    				<h3>El muchacho se tomó una selfie mientras su pareja le era infiel y luego publicó la reacción de su ahora exnovia.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_10">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/director-de-guardianes-de-la-galaxia-confiesa-la-triste-verdad-sobre-groot-50952">
					<h2>Director de "Guardianes de la Galaxia" confiesa la triste verdad sobre Groot</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/director-de-guardianes-de-la-galaxia-confiesa-la-triste-verdad-sobre-groot-50952"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/director-de-guardianes-de-la-galaxia-confiesa-la-triste-verdad-sobre-groot-50952" sharetext="Director de "Guardianes de la Galaxia" confiesa la triste verdad sobre Groot #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/director-de-guardianes-de-la-galaxia-confiesa-la-triste-verdad-sobre-groot-50952"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/director-de-guardianes-de-la-galaxia-confiesa-la-triste-verdad-sobre-groot-50952">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5a9715577411f553d721823c.jpg" class="img_def lazy" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot">
						<noscript><img src="http://cdn.canal12.com.sv/files/5a9715577411f553d721823c.jpg" class="img_def" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5a9715577411f553d721823c.jpg" class="img_small lazy" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5a9715577411f553d721823c.jpg" class="img_small" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5a9715577411f553d721823c.jpg" class="img_tiny lazy" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5a9715577411f553d721823c.jpg" class="img_tiny" alt="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot" title="Director de Guardianes de la Galaxia confiesa la triste verdad sobre Groot"></noscript>
					</div>
    				<h3>Al parecer, muchos estaban equivocados respecto a lo que ocurrió con el querido personaje en el primer film de la saga.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article></td>
		<td id="columna_3">
            <table class="bloquenotas" style="margin-top:0px !important; border:0px !important;">
                <tr>
                    <td class="botonad" style="border:0px !important; border-bottom:1px #d8d8d8 solid !important;">
            <!-- Canal9_Portada_Boton -->
<div id='div-gpt-ad-boton'>
<script type='text/javascript'>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-boton'); });
</script>
</div>
                    </td>
                </tr>
                <tr>
                    <td style="border:0px !important;"><article class="item" id="article_1_5">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/revelan-la-verdadera-edad-que-tendrian-los-simpson-si-realmente-envejecieran-51391">
					<h2>Revelan la verdadera edad que tendrían "Los Simpson" si realmente envejecieran</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/revelan-la-verdadera-edad-que-tendrian-los-simpson-si-realmente-envejecieran-51391"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/revelan-la-verdadera-edad-que-tendrian-los-simpson-si-realmente-envejecieran-51391" sharetext="Revelan la verdadera edad que tendrían "Los Simpson" si realmente envejecieran #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/revelan-la-verdadera-edad-que-tendrian-los-simpson-si-realmente-envejecieran-51391"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/revelan-la-verdadera-edad-que-tendrian-los-simpson-si-realmente-envejecieran-51391">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa68ad37411f50fa7c6fd0b.jpg" class="img_def lazy" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa68ad37411f50fa7c6fd0b.jpg" class="img_def" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa68ad37411f50fa7c6fd0b.jpg" class="img_small lazy" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa68ad37411f50fa7c6fd0b.jpg" class="img_small" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa68ad37411f50fa7c6fd0b.jpg" class="img_tiny lazy" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa68ad37411f50fa7c6fd0b.jpg" class="img_tiny" alt="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran" title="Revelan la verdadera edad que tendrían Los Simpson si realmente envejecieran"></noscript>
					</div>
    				<h3>Los fanáticos de esta exitosa serie siempre han querido saber cuántos años tendrían sus personajes y, al fin, se resolvió el misterio.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_8">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/la-fuerte-imagen-de-arnold-schwarzenegger-a-los-16-anos-que-sorprende-a-sus-fans -51388">
					<h2>La "fuerte" imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans </h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/la-fuerte-imagen-de-arnold-schwarzenegger-a-los-16-anos-que-sorprende-a-sus-fans -51388"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/la-fuerte-imagen-de-arnold-schwarzenegger-a-los-16-anos-que-sorprende-a-sus-fans -51388" sharetext="La "fuerte" imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans  #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/la-fuerte-imagen-de-arnold-schwarzenegger-a-los-16-anos-que-sorprende-a-sus-fans -51388"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/la-fuerte-imagen-de-arnold-schwarzenegger-a-los-16-anos-que-sorprende-a-sus-fans -51388">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5aa68aed7411f50fa7c6fd39.jpg" class="img_def lazy" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans ">
						<noscript><img src="http://cdn.canal12.com.sv/files/5aa68aed7411f50fa7c6fd39.jpg" class="img_def" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans "></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5aa68aed7411f50fa7c6fd39.jpg" class="img_small lazy" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans ">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5aa68aed7411f50fa7c6fd39.jpg" class="img_small" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans "></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5aa68aed7411f50fa7c6fd39.jpg" class="img_tiny lazy" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans ">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5aa68aed7411f50fa7c6fd39.jpg" class="img_tiny" alt="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans " title="La fuerte imagen de Arnold Schwarzenegger a los 16 años que sorprende a sus fans "></noscript>
					</div>
    				<h3>El actor demostró que desde su adolescencia se interesó por fortalecer y tonificar su cuerpo.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article><article class="item" id="article_1_11">
				<a class="enlace" href="http://www.canal12.com.sv/espectaculos/los-desconocidos-detalles-para-lograr-una-perfecta-ceremonia-de-los-premios-oscar-50928">
					<h2>Los desconocidos detalles para lograr una "perfecta" ceremonia de los premios Oscar</h2>
				</a>
    			<div class="fecha"></div>
				<div class="redes">
					<div class="cab">Compartir en:</div>
					<div class="share fb">
						<div class="ico fb" id="fblink" sharelink="https://www.facebook.com/sharer/sharer.php?u=http://www.canal12.com.sv/espectaculos/los-desconocidos-detalles-para-lograr-una-perfecta-ceremonia-de-los-premios-oscar-50928"></div>
					</div>
					<div class="share tw">
						<div class="ico tw" id="twlink" sharelink="http://www.canal12.com.sv/espectaculos/los-desconocidos-detalles-para-lograr-una-perfecta-ceremonia-de-los-premios-oscar-50928" sharetext="Los desconocidos detalles para lograr una "perfecta" ceremonia de los premios Oscar #ElSalvador via @#"></div>
					</div>
					<div class="share gp">
						<div class="ico gp" id="gplink" sharelink="https://plus.google.com/share?url=http://www.canal12.com.sv/espectaculos/los-desconocidos-detalles-para-lograr-una-perfecta-ceremonia-de-los-premios-oscar-50928"></div>
					</div>
				</div>
				<a href="http://www.canal12.com.sv/espectaculos/los-desconocidos-detalles-para-lograr-una-perfecta-ceremonia-de-los-premios-oscar-50928">
					<div class="imgart">
						<div class="shadowbox">
							<div class="icono foto" style="display:none"></div>
							<div class="icono video" style="display:none"></div>
						</div>
						<img data-original="http://cdn.canal12.com.sv/files/5a96d2297411f553d7217627.jpg" class="img_def lazy" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar">
						<noscript><img src="http://cdn.canal12.com.sv/files/5a96d2297411f553d7217627.jpg" class="img_def" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/316x202_5a96d2297411f553d7217627.jpg" class="img_small lazy" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar">
						<noscript><img src="http://cdn.canal12.com.sv/files/316x202_5a96d2297411f553d7217627.jpg" class="img_small" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar"></noscript>
						<img data-original="http://cdn.canal12.com.sv/files/175x112_5a96d2297411f553d7217627.jpg" class="img_tiny lazy" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar">
						<noscript><img src="http://cdn.canal12.com.sv/files/175x112_5a96d2297411f553d7217627.jpg" class="img_tiny" alt="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar" title="Los desconocidos detalles para lograr una perfecta ceremonia de los premios Oscar"></noscript>
					</div>
    				<h3>Son cientos de personas las que trabajan para que la jornada resulte lo mejor posible y sin errores.</h3>
    				<div class="frase"><span></span></div>
    			</a>
			</article></td>
                </tr>
            </table>
        </td>
	</tr>
</table></section>

<footer id="footer">
  <div class="row footer">
    <div class="mapasitio">
      <ul class="lista">
        <li><a href="" class="cab">INICIO</a></li>
        <li><a href="/envivo">En Vivo</a></li>
        <li><a href="/programas">Programas</a></li>
        <li><a href="/novelas">Novelas</a></li>
      </ul>
      <ul class="lista">
        <li><a href="/noticias/actualidad-1" class="cab">ACTUALIDAD</a></li>
        <li><a href="/noticias/nacionales-3068">Nacionales</a></li>
        <li><a href="/noticias/internacional-3069">Internacional</a></li>
        <li><a href="/noticias/sucesos-3070">Sucesos</a></li>
        <li><a href="/noticias/economia-3071">Economía</a></li>
        <li><a href="/noticias/salud-3072">Salud</a></li>
        <li><a href="/noticias/politica-3073">Política</a></li>
        <li><a href="/noticias/tecnologia-3074">Tecnología</a></li>
        <li><a href="/noticias/cultura-3075">Cultura</a></li>
        <li><a href="/noticias/reportajes-3076">Reportajes</a></li>
        <li><a href="/noticias/cocina-3077">Cocina</a></li>
        <li><a href="/noticias/variedades-3078">Variedades</a></li>
        <li><a href="/noticias/redes-sociales-3078">Redes Sociales</a></li>
      </ul>
      <ul class="lista">
        <li><a href="/noticias/deportes-3" class="cab">DEPORTES</a></li>
        <li><a href="/noticias/futbol-nacional-3064">Fútbol Nacional</a></li>
        <li><a href="/noticias/futbol-internacional-3065">Fútbol Internacional</a></li>
        <li><a href="/noticias/seleccion-nacional-3066">Selección Nacional</a></li>
        <li><a href="/noticias/mas-deportes-3067">Más Deportes</a></li>
      </ul>
      <ul class="lista">
        <li><a href="/noticias/espectaculos-2" class="cab">ESPECTACULOS</a></li>
        <li><a href="/noticias/cine-3080">Cine</a></li>
        <li><a href="/noticias/entretenimiento-3081">Entretenimiento</a></li>
        <li><a href="/noticias/musica-3082">Música</a></li>
      </ul>
    </div>
    <div class="pieiconos">
      <div class="izq"> <a href="" target="_blank" class="logo"></a>
        <div class="search">
          <input type="text" class="tbuscador">
          <div class="btnsearch">
            <div class="ico"></div>
          </div>
        </div>
        <div class="enlaces">
          <div>Derechos Reservados Red El Salvador S.A. 2015</div>
          <div> <a href="/contactenos" class="link borde">CONTÁCTENOS</a> </div>
        </div>
      </div>
      <div class="der">
        <div class="redes"> <span class="texto">Síguenos en</span>
          <ul>
            <li><a href="http://www.facebook.com/CanalDoceSV" class="fb" target="_blank"></a></li>
            <li><a href="http://www.twitter.com/Canal_12" class="tw" target="_blank"></a></li>
            <li><a href="http://plus.google.com/100912321241699444897" class="gp" target="_blank"></a></li>
            <li><a href="https://www.youtube.com/canal12sv" class="yt" target="_blank"></a></li>
          </ul>
        </div>
        <div class="grupo">
          <div class="logogrupo"></div>
          <div class="texto">Red El Salvador S.A.<br>
            El Salvador</div>
        </div>
        <div class="canales">
          <ul>
            <li class="ico atv"></li>
            <li class="ico global"></li>
            <li class="ico latele"></li>
            <li class="ico atvmas"></li>
            <li class="ico atvsur"></li>
          </ul>
        </div>
      </div>
    </div>
  </div>
</footer><script language="javascript" type="text/javascript">
$(function() {
    $("img.lazy").lazyload({
		effect : "fadeIn",
    	threshold : 200,
		failure_limit : 10
	});
});
</script>
</body>
</html>