

<!-- ////HOME/// -->

<!DOCTYPE html>
<html prefix="og: http://ogp.me/ns#" xmlns="http://www.w3.org/1999/xhtml" xml:lang="es-es" lang="es-es" dir="ltr">
<head>
	<meta name="viewport" content="width=device-width, initial-scale=1.0" />
	<meta http-equiv="X-UA-Compatible" content="IE=edge">
	  <base href="http://www.mined.gob.sv/" />
  <meta http-equiv="content-type" content="text/html; charset=utf-8" />
  <meta name="keywords" content="mined, ministerio de educación,educación,niños,escuela,paes,colección cipotes, planes de estudio" />
  <meta name="rights" content="Ministerio de Educación,Todos los derechos reservados , Gobierno de El Salvador Edificios A, Plan Maestro, Centro de Gobierno, Alameda Juan Pablo II y calle Guadalupe, San Salvador, El Salvador, América Central. Teléfonos: +(503) 2592-2000, +(503) 2592-2122, +(503) 2592-3117 Correo electrónico: educacion@mined.gob.sv Mapa de Ubicación" />
  <meta name="description" content="Ministerio de Educación El Salvador" />
  <title>Inicio</title>
  <link href="http://www.mined.gob.sv/index.php" rel="canonical" />
  <link href="/index.php?format=feed&amp;type=rss" rel="alternate" type="application/rss+xml" title="RSS 2.0" />
  <link href="/index.php?format=feed&amp;type=atom" rel="alternate" type="application/atom+xml" title="Atom 1.0" />
  <link href="/templates/protostar/favicon.ico" rel="shortcut icon" type="image/vnd.microsoft.icon" />
  <link href="http://www.mined.gob.sv/index.php/component/search/?layout=blog&amp;id=2&amp;Itemid=101&amp;format=opensearch" rel="search" title="Buscar Ministerio de Educación" type="application/opensearchdescription+xml" />
  <link rel="stylesheet" href="/components/com_k2/css/k2.css" type="text/css" />
  <link rel="stylesheet" href="/templates/protostar/css/template.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_carousel_banner/assets/css/flexisel.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_slideshowck/themes/default/css/camera.css" type="text/css" />
  <link rel="stylesheet" href="https://fonts.googleapis.com/css?family=Droid+Sans" type="text/css" />
  <link rel="stylesheet" href="http://www.mined.gob.sv/modules/mod_icemegamenu/themes/clean/css/clean_icemegamenu.css" type="text/css" />
  <link rel="stylesheet" href="http://www.mined.gob.sv/modules/mod_icemegamenu/themes/clean/css/clean_icemegamenu-reponsive.css" type="text/css" />
  <link rel="stylesheet" href="/media/jfontsize/css/jfontsize.css" type="text/css" />
  <style type="text/css">

        #mycarousel-121 {display:none;}
        .nbs-flexisel-item img { max-width:468; max-height:60;}
    #camera_wrap_100 .camera_pag_ul li img, #camera_wrap_100 .camera_thumbs_cont ul li > img {height:75px;}
#camera_wrap_100 .camera_caption {
	display: block;
	position: absolute;
}
#camera_wrap_100 .camera_caption > div {
	font-size: 12px;font-family:'Droid Sans';
}
#camera_wrap_100 .camera_caption > div div.slideshowck_description {
	font-size: 10px;
}

@media screen and (max-width: 480px) {
		.camera_caption {
			display: none !important;
		}
}
  </style>
  <script src="/media/system/js/mootools-core.js" type="text/javascript"></script>
  <script src="/media/system/js/core.js" type="text/javascript"></script>
  <script src="/media/jui/js/jquery.min.js" type="text/javascript"></script>
  <script src="/media/jui/js/jquery-noconflict.js" type="text/javascript"></script>
  <script src="/media/jui/js/jquery-migrate.min.js" type="text/javascript"></script>
  <script src="/components/com_k2/js/k2.js?v2.6.9&amp;sitepath=/" type="text/javascript"></script>
  <script src="/media/system/js/caption.js" type="text/javascript"></script>
  <script src="/media/jui/js/bootstrap.min.js" type="text/javascript"></script>
  <script src="/templates/protostar/js/template.js" type="text/javascript"></script>
  <script src="/modules/mod_carousel_banner/assets/js/jquery.noconflict.js" type="text/javascript"></script>
  <script src="/modules/mod_carousel_banner/assets/js/jquery.flexisel.js" type="text/javascript"></script>
  <script src="/modules/mod_slideshowck/assets/jquery.easing.1.3.js" type="text/javascript"></script>
  <script src="/modules/mod_slideshowck/assets/jquery.mobile.customized.min.js" type="text/javascript"></script>
  <script src="/modules/mod_slideshowck/assets/camera.min.js" type="text/javascript"></script>
  <script src="/media/jfontsize/js/jquery.jfontsize-1.0.min.js" type="text/javascript"></script>
  <script src="/media/system/js/html5fallback.js" type="text/javascript"></script>
  <script type="text/javascript">
jQuery(window).on('load',  function() {
				new JCaption('img.caption');
			});
    jQuery(window).load(function() {
        jQuery("#mycarousel-121").flexisel({

                visibleItems: 5, // $visible_items
                animationSpeed: 3000, // 1000
                autoPlay: 1, // false
                autoPlaySpeed:  1000, // 3000
                pauseOnHover: 1, // true
                enableResponsiveBreakpoints: true,
                responsiveBreakpoints: {
                    portrait: {
                        changePoint:480,
                        visibleItems: 2
                    },
                    landscape: {
                        changePoint:640,
                        visibleItems: 4
                    },
                    tablet: {
                        changePoint:768,
                        visibleItems: 1
                    }
                }
            });
        });
    
  </script>
  <script type="text/javascript">
	(function ($) {
		$().ready(function () {
			 $('body').jfontsize({
			     btnMinusClasseId: '#jfontsize-minus',
			     btnDefaultClasseId: '#jfontsize-default',
			     btnPlusClasseId: '#jfontsize-plus',
			     btnMinusMaxHits: 10,
			     btnPlusMaxHits: 10,
			     sizeChange: 1
			 });
		});
	})(jQuery)
</script>

					<style type="text/css">
		body.site
		{
			border-top: 3px solid #0088cc;
		}
		a{
			color: #0088cc;
		}
		
		
	</style>
		<!--[if lt IE 9]>
		<script src="/media/jui/js/html5.js"></script>
	<![endif]-->

</head>

<body class="site com_content view-category layout-blog no-task itemid-101">

<!--<center>
<a href="http://distancia.ues.edu.sv/" target="_blank">
<img src="/images/uonline.jpg"/>
</a>
</center>-->

<!-- Body -->
<div class="body">

<div class="container">
<!-- Header -->
<header class="header" role="banner">

<!--INICIO CONTROLES-->
<div class="row-fluid" style="border-bottom:1px solid #ccc">
	<div class="span12">
		<div class="span4"> 
			<!--		<div class="moduletable">
						<div class="search">
	<form action="/index.php" method="post" class="form-inline">
		<label for="mod-search-searchword" class="element-invisible">Buscar</label> <input name="searchword" id="mod-search-searchword" maxlength="200"  class="inputbox search-query" type="search" size="20" placeholder="Buscar" />		<input type="hidden" name="task" value="search" />
		<input type="hidden" name="option" value="com_search" />
		<input type="hidden" name="Itemid" value="101" />
	</form>
</div>
		</div>
	-->
<!---->

<script>
  (function() {
    var cx = '016356521776151587337:fgtbghisok4';
    var gcse = document.createElement('script');
    gcse.type = 'text/javascript';
    gcse.async = true;
    gcse.src = 'https://cse.google.com/cse.js?cx=' + cx;
    var s = document.getElementsByTagName('script')[0];
    s.parentNode.insertBefore(gcse, s);
  })();
</script>
<gcse:search></gcse:search>

<!---->
		</div>
		<div class="span2"> 		<div class="moduletable social">
						<!-- BEGIN: Custom advanced (www.pluginaria.com) -->
<a name="participacion" href="http://twitter.com/MINEDelsalvador"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-twitter fa-stack-1x fa-inverse"></i>
          </span>
</a> 
<a name="participacion" href="https://www.facebook.com/MINEDelsalvador"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-facebook fa-stack-1x fa-inverse"></i>
          </span>
</a>
<a name="participacion" href="https://www.youtube.com/channel/UC7JZ4j5-dQX6j8BgaASOP_Q"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-youtube fa-stack-1x fa-inverse"></i>
          </span>
</a> 
    <!-- END: Custom advanced (www.pluginaria.com) -->
		</div>
	</div>
		<div class="span1">  </div>
        	<div class="span2">		<div class="moduletable">
						<div class="jfontsize">
	<a class="jfontsize-button" id="jfontsize-minus">A-</a>
	<a class="jfontsize-button" id="jfontsize-default">A</a>
	<a class="jfontsize-button" id="jfontsize-plus">A+</a>
</div>		</div>
	</div>
		
		<div class="span3" style="background: #004f7d;"><a href="http://publica.gobiernoabierto.gob.sv/institutions/ministerio-de-educacion" target="_blank"><img src='/images/ptransparencia.jpg'></a></div>
	</div>  
</div> 
<!--FIN CONTROLES-->   

<!-- ///// FRASE Y LOGO DEL MINED /// -->
    <div class="header-inner clearfix">
        <a class="brand pull-left span9" href="/">
				<h1 style="color:#16668f!important; font-size:35px">Ministerio de Educaci&oacute;n<br><small>Rep&uacute;blica de El Salvador</small></h1>
                        </a>
	<div class="span3 logo-mined"><img src="/images/alfa2018.jpg" alt="Ministerio de Educaci�n" ></div>

					
    </div>
    
		<div style="padding-left:20px;">
			
        </div>

</header><!-- FIN HEADER  -->
			
<!-- ///// MENU PRINCIPAL /// -->
			<div class="row-fluid menu">
			    <span class="hidden-desktop txt-hidden">MENU PRINCIPAL</span>
				<div class="span12 menu">
				    <div class="icemegamenu"><div class="ice-megamenu-toggle"><a data-toggle="collapse" data-target=".nav-collapse">Menu</a></div><div class="nav-collapse icemegamenu collapse  "><ul id="icemegamenu" class="meganizr mzr-slide mzr-responsive"><li id="iceMenu_101" class="iceMenuLiLevel_1 active"><a href="http://www.mined.gob.sv/" class="icemega_active iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Inicio</span></a></li><li id="iceMenu_156" class="iceMenuLiLevel_1 mzr-drop parent"><a href="#" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Institución</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_175" class="iceMenuLiLevel_2"><a href="/index.php/institucion/estructura-organizativa" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Estructura Organizativa</span></a></li><li id="iceMenu_183" class="iceMenuLiLevel_2"><a href="/index.php/institucion/marco-legal" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Marco Legal</span></a></li><li id="iceMenu_181" class="iceMenuLiLevel_2"><a href="/index.php/institucion/filosofia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Filosofía</span></a></li><li id="iceMenu_184" class="iceMenuLiLevel_2"><a href="/index.php/institucion/autoridades" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Autoridades</span></a></li><li id="iceMenu_178" class="iceMenuLiLevel_2"><a href="/index.php/institucion/transparencia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Transparencia</span></a></li><li id="iceMenu_186" class="iceMenuLiLevel_2"><a href="https://webmail.mined.gob.sv/owa/" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Área Institucional</span></a></li></ul></div></li></ul></li><li id="iceMenu_127" class="iceMenuLiLevel_1 mzr-drop parent"><a href="/index.php/servicios" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Servicios</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_332" class="iceMenuLiLevel_2"><a href="http://www.mined.gob.sv/index.php/descargas/category/942-servicios" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Colegios Privados</span></a></li><li id="iceMenu_188" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/406-división-de-legalización-de-centros-educativos" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">División de legalización de centros educativos </span></a></li><li id="iceMenu_189" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/407-atención-a-necesidades-educativas-especiales" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Atención a necesidades educativas especiales </span></a></li><li id="iceMenu_190" class="iceMenuLiLevel_2"><a href="/index.php/servicios/educacion-superior" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Educación Superior </span></a></li><li id="iceMenu_191" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/409-registro-e-incorporaciones" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Registro e Incorporaciones</span></a></li><li id="iceMenu_192" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/410-asesoría-jurídica" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Asesoría Jurídica</span></a></li><li id="iceMenu_193" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/411-división-de-estudios" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">División de Estudios </span></a></li><li id="iceMenu_194" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/412-división-de-formación-docente" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">División de Formación Docente </span></a></li><li id="iceMenu_196" class="iceMenuLiLevel_2"><a href="/index.php/servicios/itemlist/category/483-educación-media" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Educación Media</span></a></li><li id="iceMenu_197" class="iceMenuLiLevel_2"><a href="/index.php/servicios/en-linea" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">En línea</span></a></li><li id="iceMenu_283" class="iceMenuLiLevel_2"><a href="/index.php/servicios/sistema-georeferencia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Sistema Georeferencia</span></a></li><li id="iceMenu_293" class="iceMenuLiLevel_2"><a href="/index.php/servicios/busqueda-de-planes" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Busqueda de planes de estudio y universidades autorizadas</span></a></li></ul></div></li></ul></li><li id="iceMenu_128" class="iceMenuLiLevel_1 mzr-drop parent"><a href="/index.php/noticias" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Noticias</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_204" class="iceMenuLiLevel_2"><a href="/index.php/noticias/historial-de-noticias" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Historial de Noticias</span></a></li><li id="iceMenu_206" class="iceMenuLiLevel_2"><a href="/index.php/noticias/avisos" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Avisos</span></a></li><li id="iceMenu_207" class="iceMenuLiLevel_2"><a href="https://www.youtube.com/channel/UC7JZ4j5-dQX6j8BgaASOP_Q" target="_blank" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Multimedia</span></a></li><li id="iceMenu_337" class="iceMenuLiLevel_2"><a href="/index.php/noticias/alfabetizacion" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Alfabetización</span></a></li></ul></div></li></ul></li><li id="iceMenu_141" class="iceMenuLiLevel_1"><a href="/index.php/descargas" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Descargas</span></a></li><li id="iceMenu_157" class="iceMenuLiLevel_1 mzr-drop parent"><a href="/index.php/programas-educativos" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programas Educativos</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_312" class="iceMenuLiLevel_2 mzr-drop parent"><a href="#" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Ciencia y Tecnología</span></a><ul class="icesubMenu icemodules sub_level_2" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_199" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/aeds.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Atención a Estudiantes con Desempeño Sobresaliente</span></a></li><li id="iceMenu_311" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/ppc.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa Presidencial "Una Niña, Un Niño, Una Computadora"</span></a></li><li id="iceMenu_313" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/ensanche.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa Ensanche de las Tecnologías de La Información y Comunicación y su Uso Responsable (Ensanche)</span></a></li><li id="iceMenu_314" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/cyma.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Sub Programa “Hacia La Cyma”</span></a></li><li id="iceMenu_315" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/psp.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa Seamos Productivos</span></a></li><li id="iceMenu_316" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/snetp.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Fortalecimiento del Sistema de Formación Técnico Profesional</span></a></li><li id="iceMenu_317" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/pse.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Subrograma Sigamos Estudiando</span></a></li><li id="iceMenu_319" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/sbg.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Subprograma Becas GOES</span></a></li><li id="iceMenu_320" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/sistema-de-seguimiento-a-la-calidad-educativa.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Subprograma Sistema de Seguimiento a la Calidad</span></a></li><li id="iceMenu_321" class="iceMenuLiLevel_3"><a href="http://www.cienciaytecnologia.edu.sv/programas/pcc.html" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa Creando Conocimiento</span></a></li></ul></div></li></ul></li><li id="iceMenu_202" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/eitp" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Escuela Inclusiva de Tiempo Pleno</span></a></li><li id="iceMenu_203" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/educacion-superior" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Educación Superior</span></a></li><li id="iceMenu_282" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/formacion-docente" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Formación docente</span></a></li><li id="iceMenu_288" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/ajedrez-educativo" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Ajedrez Educativo</span></a></li><li id="iceMenu_289" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/dnge" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Gestión Educativa</span></a></li><li id="iceMenu_304" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/unidad-de-genero" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Política de Género</span></a></li><li id="iceMenu_308" class="iceMenuLiLevel_2"><a href="http://distancia.ues.edu.sv/" target="_blank" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Universidad en Línea</span></a></li><li id="iceMenu_309" class="iceMenuLiLevel_2"><a href="/index.php/programas-sociales/item/7913-sub-programa-vaso-de-leche" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Vaso de Leche</span></a></li><li id="iceMenu_310" class="iceMenuLiLevel_2"><a href="/index.php/programas-sociales/item/5480-programa-de-alimentacion-y-salud-escolar" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa de Alimentación y Salud Escolar</span></a></li><li id="iceMenu_198" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/paquete-escolar" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Paquete Escolar</span></a></li><li id="iceMenu_200" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/programa-de-alfabetizacion" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa de Alfabetización</span></a></li><li id="iceMenu_326" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/maesre" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Mejoramiento de los Ambientes Escolares y Recursos Educativos</span></a></li><li id="iceMenu_327" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/educacion-ambiental-gestion-de-riesgos-y-cambio-climatico" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Educación Ambiental, Gestión de Riesgos y Cambio Climático</span></a></li><li id="iceMenu_328" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/programa-de-inmersion-lingueistica-temprana-cuna-nahuat" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Programa de Inmersión Lingüística Temprana, Cuna Náhuat</span></a></li><li id="iceMenu_329" class="iceMenuLiLevel_2"><a href="/index.php/programas-educativos/esmate" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Proyecto de Mejoramiento de Aprendizajes en Matemática en Educación Básica y Educación Media (ESMATE)</span></a></li></ul></div></li></ul></li><li id="iceMenu_158" class="iceMenuLiLevel_1 mzr-drop parent"><a href="#" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Contáctenos</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_208" class="iceMenuLiLevel_2"><a href="/index.php/contactenos/buzon-de-sugerencias" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Buzón de Sugerencias</span></a></li><li id="iceMenu_209" class="iceMenuLiLevel_2"><a href="#participacion" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Participación Ciudadana</span></a></li><li id="iceMenu_210" class="iceMenuLiLevel_2"><a href="/index.php/contactenos/esquema-oficinas-centrales" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Esquema de Oficinas Centrales</span></a></li><li id="iceMenu_211" class="iceMenuLiLevel_2"><a href="/index.php/contactenos/oficinas-departamentales" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Oficinas Departamentales</span></a></li><li id="iceMenu_212" class="iceMenuLiLevel_2"><a href="/index.php/contactenos/direcorio-ce" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Directorio de Centros Educativos</span></a></li></ul></div></li></ul></li><li id="iceMenu_213" class="iceMenuLiLevel_1 mzr-drop parent"><a href="#" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Ayuda</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_214" class="iceMenuLiLevel_2"><a href="/index.php/2015-05-13-22-38-34/preguntas-frecuentes" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Preguntas Frecuentes</span></a></li><li id="iceMenu_215" class="iceMenuLiLevel_2"><a href="/index.php/2015-05-13-22-38-34/buscador" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Buscador</span></a></li><li id="iceMenu_216" class="iceMenuLiLevel_2"><a href="/index.php/2015-05-13-22-38-34/politica-uso-de-documentos-y-recursos-publicados" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Política Uso de Documentos y Recursos Publicados</span></a></li><li id="iceMenu_270" class="iceMenuLiLevel_2"><a href="/index.php/2015-05-13-22-38-34/carta-de-derechos" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Carta de derechos</span></a></li><li id="iceMenu_271" class="iceMenuLiLevel_2"><a href="/index.php/2015-05-13-22-38-34/politica-de-seguridad" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Politica de seguridad y privacidad de datos</span></a></li></ul></div></li></ul></li><li id="iceMenu_266" class="iceMenuLiLevel_1 mzr-drop parent"><a href="#" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Area Interna</span></a><ul class="icesubMenu  sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_267" class="iceMenuLiLevel_2"><a href="http://sistemas.mined.gob.sv/sae/login.do;jsessionid=4F49FA89C19F204AE873A37C1C8386FC" target="_blank" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">SAE</span></a></li><li id="iceMenu_268" class="iceMenuLiLevel_2"><a href="http://intranet.mined.gob.sv" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Intranet</span></a></li><li id="iceMenu_269" class="iceMenuLiLevel_2"><a href="https://webmail.mined.gob.sv/owa/auth/logon.aspx?url=https://webmail.mined.gob.sv/owa/&amp;reason=0" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Correo Institucional</span></a></li><li id="iceMenu_159" class="iceMenuLiLevel_2"><a href="/index.php/area-interna/funcionarios" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Funcionarios</span></a></li><li id="iceMenu_295" class="iceMenuLiLevel_2"><a href="/index.php/area-interna/manual-de-servicios-y-prestaciones" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Manual de servicios y prestaciones</span></a></li><li id="iceMenu_323" class="iceMenuLiLevel_2"><a href="/descarga/Procedimiento Administrativo MINED.pdf" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Procedimiento Administrativo MINED</span></a></li></ul></div></li></ul></li><li id="iceMenu_286" class="iceMenuLiLevel_1 mzr-drop parent"><a href="/index.php/paes-cat" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">PAES</span></a><ul class="icesubMenu icemodules sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_335" class="iceMenuLiLevel_2"><a href="/index.php/paes-cat/actualizacion-em" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Actualización de datos educación media</span></a></li></ul></div></li></ul></li></ul></div></div>


<script type="text/javascript">
	jQuery(document).ready(function(){
		var browser_width1 = jQuery(window).width();
		jQuery("#icemegamenu").find(".icesubMenu").each(function(index){
			var offset1 = jQuery(this).offset();
			var xwidth1 = offset1.left + jQuery(this).width();
			if(xwidth1 >= browser_width1){
				jQuery(this).addClass("ice_righttoleft");
			}
		});
		
	})
	jQuery(window).resize(function() {
		var browser_width = jQuery(window).width();
		jQuery("#icemegamenu").find(".icesubMenu").removeClass("ice_righttoleft");
		jQuery("#icemegamenu").find(".icesubMenu").each(function(index){
			var offset = jQuery(this).offset();
			var xwidth = offset.left + jQuery(this).width();
			
			if(xwidth >= browser_width){
				jQuery(this).addClass("ice_righttoleft");
			}
		});
	});
</script>
				</div>
			</div>
	
<!-- ///// SLIDE /// -->
			<div class="row-fluid">
				<div class="span12">
							<div class="moduletable">
						
		<!--[if lte IE 7]>
		<link href="/modules/mod_slideshowck/themes/default/css/camera_ie.css" rel="stylesheet" type="text/css" />
		<![endif]-->
		<!--[if IE 8]>
		<link href="/modules/mod_slideshowck/themes/default/css/camera_ie8.css" rel="stylesheet" type="text/css" />
		<![endif]--><script type="text/javascript"> <!--
       jQuery(function(){
        jQuery('#camera_wrap_100').camera({
                height: '345px',
                minHeight: '',
                pauseOnClick: false,
                hover: 1,
                fx: 'simpleFade',
                loader: 'none',
                pagination: 0,
                thumbnails: 0,
                thumbheight: 75,
                thumbwidth: 100,
                time: 7000,
                transPeriod: 1500,
                alignment: 'bottomLeft',
                autoAdvance: 1,
                mobileAutoAdvance: 1,
                portrait: 0,
                barDirection: 'leftToRight',
                imagePath: '/modules/mod_slideshowck/images/',
                lightbox: 'mediaboxck',
                fullpage: 0,
				mobileimageresolution: '640',
                navigationHover: true,
				mobileNavHover: true,
				navigation: true,
				playPause: true,
                barPosition: 'bottom',
				container: ''
        });
}); //--> </script><!-- debut Slideshow CK -->
<div class="slideshowck camera_wrap camera_black_skin" id="camera_wrap_100">
			<div data-rel="lightbox" data-thumb="/images/th/ASFM_th.jpg" data-src="/images/ASFM.jpg" data-link="http://www.mined.gob.sv/index.php/noticias/item/9325-buscan-alfabetizar-a-695-personas-en-san-francisco-menendez" data-target="lightbox" data-alignment="topCenter">
							<div class="camera_caption fadeIn">
					<div class="camera_caption_title">
						Buscan alfabetizar a 695 personas en San Francisco Menéndez											</div>
					<div class="camera_caption_desc">
																	</div>
				</div>
					</div>
		<div data-rel="lightbox" data-thumb="/images/th/JTalen_th.jpg" data-src="/images/JTalen.jpg" data-link="http://www.mined.gob.sv/index.php/noticias/item/9324-programa-jovenes-talento-realiza-olimpiada-salvadorena-de-informatica" data-target="lightbox" data-alignment="center">
							<div class="camera_caption fadeIn">
					<div class="camera_caption_title">
						Programa Jóvenes Talento realiza Olimpiada Salvadoreña de Informática											</div>
					<div class="camera_caption_desc">
																	</div>
				</div>
					</div>
		<div data-rel="lightbox" data-thumb="/images/th/Alca_th.jpg" data-src="/images/Alca.jpg" data-link="http://www.mined.gob.sv/index.php/noticias/item/9323-mined-alfabetizara-a-15-688-personas-en-cabanas" data-target="lightbox" data-alignment="topCenter">
							<div class="camera_caption fadeIn">
					<div class="camera_caption_title">
						MINED alfabetizará a 15,688 personas en Cabañas											</div>
					<div class="camera_caption_desc">
																	</div>
				</div>
					</div>
		<div data-rel="lightbox" data-thumb="/images/th/BJ_th.jpg" data-src="/images/BJ.jpg" data-link="http://www.mined.gob.sv/index.php/noticias/item/9322-estudiante-del-programa-de-jovenes-talento-obtiene-beca-para-estudiar-en-japon" data-target="lightbox" data-alignment="center">
							<div class="camera_caption fadeIn">
					<div class="camera_caption_title">
						Estudiante del Programa de Jóvenes Talento obtiene beca para estudiar en Japón											</div>
					<div class="camera_caption_desc">
																	</div>
				</div>
					</div>
		<div data-rel="lightbox" data-thumb="/images/th/JT10_th.jpg" data-src="/images/JT10.jpg" data-link="http://www.mined.gob.sv/index.php/noticias/item/9321-dos-estudiantes-del-programa-jovenes-talento-son-aceptados-en-el-instituto-tecnologico-de-massachusetts" data-target="lightbox" data-alignment="center">
							<div class="camera_caption fadeIn">
					<div class="camera_caption_title">
						Dos estudiantes del Programa Jóvenes Talento son aceptados en el Instituto Tecnológico de Massachusetts											</div>
					<div class="camera_caption_desc">
																	</div>
				</div>
					</div>
</div>
<div style="clear:both;"></div>
<!-- fin Slideshow CK -->
		</div>
	
				</div>
			</div>


<!--  /// PROGRAMAS MINED /// -->

    <div class="row-fluid">
                <div class="span12 programa nav nav-stacked">
            <!-- BEGIN: Custom advanced (www.pluginaria.com) -->
<ul class="programas">
<li><a class= "btn-program" href="http://www.cienciaytecnologia.edu.sv">Ciencia y Tecnología</a></li>
<li><a class= "btn-program" href="/index.php/programas-educativos/formacion-docente">Formación Docente</a></li>
<li><a class= "btn-program" href="/index.php/programas-sociales">Programas Sociales</a></li>
<li><a class= "btn-program" href="/index.php/programas-educativos/programa-de-alfabetizacion">Programa Alfabetización </a></li>
<li><a class= "btn-program" href="/index.php/programas-educativos/item/3-educacion-inicial-y-desarrollo-integral-para-la-primera-infancia">Programa Primera Infancia</a></li>
<li><a class= "btn-program btn-nino" href="http://www.cienciaytecnologia.edu.sv/programas/ppc.html"> Una Niña, Un Niño <br/> Una Computadora</a></li>
<li><a class= "btn-program" href="/index.php/programas-educativos/educacion-superior">Educación Superior</a></li>
<li><a class= "btn-program" href="http://distancia.ues.edu.sv/" target="_blank">Universidad en Línea </a></li>

</ul><!-- END: Custom advanced (www.pluginaria.com) -->

        </div>
				
    </div>
<!-- End  Program MINED -->
           
            <div class="row-fluid">
                <div class="span12">
                   <div class="row-fluid">


 


                    <div class="span4">
                      <div class="row-fluid">
                    
                          <div class="span3">
                               <span class="fa-stack fa-3x">
                                  <i class="fa fa-circle fa-stack-2x orange"></i>
                                  <i class="fa fa-file-o fa-stack-1x fa-inverse"></i>
                                </span>
                            </div>
                     
                      <div class="span9"><a class="plan" href="/index.php/descargas/category/740-plan-social-educativo"> Plan Social Educativo</a>
                        
                        <p style="text-align:justify">
El desarrollo del mundo actual y futuro exige una reflexi&oacute;n sobre lo que deben se las relaciones entre el conocimiento y la familia en la sociedad, para que los esfuerzos y la responsabilidad del individuo en una realidad que cambia puedan se valorados ...

</p></div>
                       
                      </div>
                    </div>

                      <div class="span4">
                       <div class="row-fluid">
                           <div class="span3">
                               <span class="fa-stack fa-3x">
                                  <i class="fa fa-circle fa-stack-2x orange"></i>
                                  <i class="fa fa-file-text fa-stack-1x fa-inverse"></i>
                                </span>
                            </div>
                           <div class="span9"><a class="plan" href="/index.php/descargas/send/716-institucional/6247-plan-nacional-de-educacion-en-funcion-de-la-nacion">Plan Nacional de Educaci&oacute;n en funci&oacute;n de la Naci&oacute;n</a>
                               <p style="text-align:justify">
El Plan Nacional de Educaci&oacute;n en Funci&oacute;n de la Naci&oacute;n propone una serie de apuestas estrat&eacute;gicas que despliegan la ruta se&ntilde;alada por el Plan Quinquenal de Desarrollo 2014-2019... 
</p></div>
                     </div>
                    </div>
<div class="span4">
                      <div class="row-fluid">
                    
                          <div class="span3">
                               <span class="fa-stack fa-3x">
                                  <i class="fa fa-circle fa-stack-2x orange"></i>
                                  <i class="fa fa-file fa-stack-1x fa-inverse"></i>
                                </span>
                            </div>
                     
                      <div class="span9"><a class="plan" href="/jdownloads/Institucional/Plan_El_Salvador_Educado.compressed.pdf"> Plan El Salvador Educado</a>
<p style="text-align:justify">                        
Este plan educativo constituye para el Consejo Nacional de Educaci&oacute;n (CONED), una de las trascendentales apuestas que los diferentes sectores sociales del pa&iacute;s impulsar&aacute;n en la presente d&eacute;cada y est&aacute; orientado a establecer el rumbo de la pol&iacute;tica educativa de El Salvador.                        <p style="text-align:justify">
</p></div>
                       
                      </div>
                    </div>
                </div>    
                  
                </div>
                            </div>

<div class="row-fluid">
	<a href="http://www.cienciaytecnologia.edu.sv/viceministerio/datos-estadisticos-de-los-programas/dts-lmp.html" target="_blank"><img src="/images/datos-mined.jpg"/></a>
</div>


			<div class="row-fluid">
				<!-- /// Avisos /// -->
				<div class="span4">
							<div class="moduletable event">
							<h3>Avisos</h3>
						
<div id="k2ModuleBox94" class="k2ItemsBlock  event">

	
	  <ul>
        <li class="even">

      <!-- Plugins: BeforeDisplay -->
      
      <!-- K2 Plugins: K2BeforeDisplay -->
      
      

 


<!-- FECHA DE CREACION -->
     <span class="moduleItemDateCreated">Lunes, 12 Marzo 2018</span>
      <!---->
<br/>
            <a class="moduleItemTitle" href="/index.php/noticias/avisos/item/9309-taller-matematica">Invitación a taller de matemática</a>
      
      
      <!-- Plugins: AfterDisplayTitle -->
      
      <!-- K2 Plugins: K2AfterDisplayTitle -->
      
      <!-- Plugins: BeforeDisplayContent -->
      
      <!-- K2 Plugins: K2BeforeDisplayContent -->
      
      
     

      <div class="clr"></div>

      
      <div class="clr"></div>

      <!-- Plugins: AfterDisplayContent -->
      
      <!-- K2 Plugins: K2AfterDisplayContent -->
      
      

      
      
      
			
			

			
      <!-- Plugins: AfterDisplay -->
      
      <!-- K2 Plugins: K2AfterDisplay -->
      
      <div class="clr"></div>
    </li>
        <li class="odd">

      <!-- Plugins: BeforeDisplay -->
      
      <!-- K2 Plugins: K2BeforeDisplay -->
      
      

 


<!-- FECHA DE CREACION -->
     <span class="moduleItemDateCreated">Miércoles, 07 Marzo 2018</span>
      <!---->
<br/>
            <a class="moduleItemTitle" href="/index.php/noticias/avisos/item/9303-guia-para-tiendas-y-cafetines-escolares">Guía para tiendas y cafetines escolares</a>
      
      
      <!-- Plugins: AfterDisplayTitle -->
      
      <!-- K2 Plugins: K2AfterDisplayTitle -->
      
      <!-- Plugins: BeforeDisplayContent -->
      
      <!-- K2 Plugins: K2BeforeDisplayContent -->
      
      
     

      <div class="clr"></div>

      
      <div class="clr"></div>

      <!-- Plugins: AfterDisplayContent -->
      
      <!-- K2 Plugins: K2AfterDisplayContent -->
      
      

      
      
      
			
			

			
      <!-- Plugins: AfterDisplay -->
      
      <!-- K2 Plugins: K2AfterDisplay -->
      
      <div class="clr"></div>
    </li>
        <li class="even">

      <!-- Plugins: BeforeDisplay -->
      
      <!-- K2 Plugins: K2BeforeDisplay -->
      
      

 


<!-- FECHA DE CREACION -->
     <span class="moduleItemDateCreated">Martes, 06 Marzo 2018</span>
      <!---->
<br/>
            <a class="moduleItemTitle" href="/index.php/noticias/avisos/item/9300-circular-no-3-2018-referente-a-actividades-para-conmemorar-8-de-marzo">Circular No. 3/2018 referente a actividades para conmemorar 8 de marzo</a>
      
      
      <!-- Plugins: AfterDisplayTitle -->
      
      <!-- K2 Plugins: K2AfterDisplayTitle -->
      
      <!-- Plugins: BeforeDisplayContent -->
      
      <!-- K2 Plugins: K2BeforeDisplayContent -->
      
      
     

      <div class="clr"></div>

      
      <div class="clr"></div>

      <!-- Plugins: AfterDisplayContent -->
      
      <!-- K2 Plugins: K2AfterDisplayContent -->
      
      

      
      
      
			
			

			
      <!-- Plugins: AfterDisplay -->
      
      <!-- K2 Plugins: K2AfterDisplay -->
      
      <div class="clr"></div>
    </li>
        <li class="odd">

      <!-- Plugins: BeforeDisplay -->
      
      <!-- K2 Plugins: K2BeforeDisplay -->
      
      

 


<!-- FECHA DE CREACION -->
     <span class="moduleItemDateCreated">Jueves, 01 Marzo 2018</span>
      <!---->
<br/>
            <a class="moduleItemTitle" href="/index.php/noticias/avisos/item/9294-instituciones-educativas-que-serviran-como-centros-de-votacion">Instituciones educativas que servirán como centros de votación</a>
      
      
      <!-- Plugins: AfterDisplayTitle -->
      
      <!-- K2 Plugins: K2AfterDisplayTitle -->
      
      <!-- Plugins: BeforeDisplayContent -->
      
      <!-- K2 Plugins: K2BeforeDisplayContent -->
      
      
     

      <div class="clr"></div>

      
      <div class="clr"></div>

      <!-- Plugins: AfterDisplayContent -->
      
      <!-- K2 Plugins: K2AfterDisplayContent -->
      
      

      
      
      
			
			

			
      <!-- Plugins: AfterDisplay -->
      
      <!-- K2 Plugins: K2AfterDisplay -->
      
      <div class="clr"></div>
    </li>
        <li class="even lastItem">

      <!-- Plugins: BeforeDisplay -->
      
      <!-- K2 Plugins: K2BeforeDisplay -->
      
      

 


<!-- FECHA DE CREACION -->
     <span class="moduleItemDateCreated">Miércoles, 28 Febrero 2018</span>
      <!---->
<br/>
            <a class="moduleItemTitle" href="/index.php/noticias/avisos/item/9289-estudiantes-convocados-a-la-segunda-fase-de-la-xi-olimpiada-salvadorena-de-fisica">Estudiantes convocados a la segunda fase de la XI Olimpiada Salvadoreña de Física</a>
      
      
      <!-- Plugins: AfterDisplayTitle -->
      
      <!-- K2 Plugins: K2AfterDisplayTitle -->
      
      <!-- Plugins: BeforeDisplayContent -->
      
      <!-- K2 Plugins: K2BeforeDisplayContent -->
      
      
     

      <div class="clr"></div>

      
      <div class="clr"></div>

      <!-- Plugins: AfterDisplayContent -->
      
      <!-- K2 Plugins: K2AfterDisplayContent -->
      
      

      
      
      
			
			

			
      <!-- Plugins: AfterDisplay -->
      
      <!-- K2 Plugins: K2AfterDisplay -->
      
      <div class="clr"></div>
    </li>
        <li class="clearList"></li>
  </ul>
  
	
	
</div>
		</div>
	
				</div>
				
				<!-- /// Multimedia /// -->
				<div class="span4">

							<div class="moduletable">
						<style>
.headerm{ height:25px;/*background-color:#d75e01;*/ color:#d75e01/*; padding-left:8px*/;padding-right:15px; padding-bottom:10px;}
.video{ float:left}
.lista{  width: 40%;float:left; /*margin-top:10px */  padding-left: 25px;}
.mm { /*background-color:#d75e01; color:#fff*/ border-bottom:#900 solid 2px;}
.mm ,.ad ,.gl { float:left; /*padding-left:10px;*/ padding-right:10px; text-transform:uppercase/*; height:35px*/ ; /*padding-top:5px*/}
.ad{ background-color:#FFF; color:#d75e01 }
.lista ul {list-style:none; padding:0; margin:0}
.lista ul li {list-style:none; padding:0; margin:0; padding-bottom: 4px;}
.lista ul li a{ text-decoration:none}
.multimedia { width:100%}
.fecham{color:#819f38; font-size:11px;}
.hitsm{color:#819f38; font-size:11px; }
</style>
<div class="multimedia">
	<div><h3>MULTIMEDIA</h3></div><div class="headerm"> <div class="mm"><a href="/index.php/noticias/multimedia" class="mm">Videos</a></div></div>
        
	<div class="video">
  
<!--<iframe width="350" height="230" src="https://www.youtube.com/embed/a5gVB3R1THA " frameborder="0" allowfullscreen></iframe> -->
<a href="https://www.youtube.com/channel/UC7JZ4j5-dQX6j8BgaASOP_Q" target="_blank"><img src="/img/youtubeMined.jpg"/></a>
<!--<iframe width="350" height="230" src="/" frameborder="0" allowfullscreen></iframe>-->

	<!--<iframe width="350" height="230" src="https://www.youtube.com/embed/Zv6td-9d9DY" frameborder="0" allowfullscreen></iframe>-->

        
    </div>
	<div class="lista" >
    
        <div style="clear:both"></div>
	<ul>
    
        </ul>
    
    </div>
    
</div>
<div style="clear:both"></div>




		</div>
	
					
				</div>
                               <div class="span4">
							<div class="moduletable event">
							<h3>De Interés</h3>
						

<div class="custom event"  >
	<center><a href="/index.php/noticias/alfabetizacion"><img src="/images/alf2018.jpg" alt="" /></a></center></div>
		</div>
	
				</div>

				
			</div>

<!--div separacion-->
<br>
<div style="height:10px;background: url('/templates/protostar/images/line-below.png')  repeat-x; /*padding-top:10px; padding-bottom:5px*/"></div>

<!--Linea 1-->
<div class="row-fluid" style="">
    <div class="span3 bt">
        <a href="/index.php/estadisticas-educativas"><img src="/images/AD.png"></a>
        

    </div>
    <div class="span3 bt"> 
        <a href="/index.php/licitaciones"><img src="/images/AB.png"></a>
    </div>
    <div class="span3 bt">

<a href="http://www.cienciaytecnologia.edu.sv/programas/sbg.html"><img src="/images/AC.png" width="100%"></a>
    </div>
<div class="span3 bt"> 
        <a href="http://distancia.ues.edu.sv/"><img src="/images/AG.png"></a>
    </div>  
<div style="clear:both"></div>
        <!--<div style="height:10px;background: url('/templates/protostar/images/line-below.png')  repeat-x; /*padding-top:10px; padding-bottom:5px*/"></div>-->
</div>

<!--Linea 4-->

<div class="row-fluid" style="">
    <div class="span3 bt">
        <a href="/index.php/esmate"><img src="/images/AE.png" alt="" /></a>

    </div>
    <div class="span3 bt"> 
        <a href="/index.php/component/k2/item/8594" target="_blank" rel="alternate"><img src="/images/AA.png" alt="Programas Moral y C�vica" width="299" height="211" /></a>    </div>
    <div class="span3 bt">
        <a href="/index.php/descargas/send/716-institucional/6422-libro-mas-alla-de-las-letras" target="_blank" rel="alternate"><img src="/images/AF.png" alt="Programas Moral y C�vica" /></a>
    </div>
<div class="span3 bt">
        <a href="http://www.mined.gob.sv/descarga/CALENDARIO_22_ENERO_2018_PRELIMINAR.pdf" target="_blank" rel="alternate"><img src="/images/AH.png" alt="Programas Moral y C�vica" /></a>
    </div>

   
<div style="clear:both"></div>
    
        <div style="height:10px;background: url('/templates/protostar/images/line-below.png')  repeat-x; /*padding-top:10px; padding-bottom:5px*/"></div>
    
</div>

<div class="row-fluid">
	<div class="span12">
				<div class="moduletable">
						
	<ul id="mycarousel-121">
		
		
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/10" target="_blank" title="Memoria de labores">
								
						
						

						<img
							src="http://www.mined.gob.sv//images/memoria_tmb.jpg"
							alt="Memoria de labores" title="" 
						/>	

					</a>						
			</li>
										
			
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/1" target="_blank" title="Educación Intergral">
								
						
						

						<img
							src="http://www.mined.gob.sv/images/banners/educacion2.jpg"
							alt="Educación Integral" title="" 
						/>	

					</a>						
			</li>
										
			
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/17" target="_blank" title="paz">
								
						
						

						<img
							src="http://www.mined.gob.sv//images/cultura.gif"
							alt="paz" title="" 
						/>	

					</a>						
			</li>
										
			
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/13" target="_blank" title="Ajedres">
								
						
						

						<img
							src="http://www.mined.gob.sv/images/banners/ajedrez.jpg"
							alt="Ajedres" title="" 
						/>	

					</a>						
			</li>
										
			
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/16" target="_blank" title="coned">
								
						
						

						<img
							src="http://www.mined.gob.sv//images/coned_tmb.jpg"
							alt="coned" title="" 
						/>	

					</a>						
			</li>
										
			
			<li>

									
						
							<!-- open in a new window -->
							<a href="/index.php/component/banners/click/18" target="_blank" title="PESS">
								
						
						

						<img
							src="http://www.mined.gob.sv//images/pess_tmb.jpg"
							alt="PESS" title="" 
						/>	

					</a>						
			</li>
										
						
	</ul><!-- end wrapper -->		</div>
	
	<div class="row-fluid">
<div class="span12">
		<!--<a href="http://www.presidencia.gob.sv/informes-de-gabinetes/"><img src="/images/polvora.jpg"/></a>-->
	</div>
	<!--<div class="span4">
		<a href="/downloads/convocatoria-9CTNI-espanol.pdf" target="_blank"><img src="/images/talento.jpg"/></a>
	</div>-->
</div>
<!--<img src="/images/polvora.jpg"/>
<br><br>-->
<div style="background-color:#02224b; color:#FFF;padding:15px;font-weight:bold;text-align:center;font-size:26px;">PROYECTOS DE GOBIERNO</div>
			<div class="proyectosGob">
		      	<a href="http://www.presidencia.gob.sv/wp-content/uploads/2015/01/Plan-Quinquenal-de-Desarrollo.pdf" target="_blank" >
				<img src="/images/proyectos_de_gobierno/1.jpg" width="220px"></a>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;
		     	<a href="http://www.presidencia.gob.sv/directorio/"><img src="/images/proyectos_de_gobierno/2.jpg" width="200px" target="_blank"></a>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;
		     	<a href="http://tves.sv/"><img src="/images/proyectos_de_gobierno/3.jpg" width="200px" target="_blank"></a>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;
		     	<a href="http://rnes.sv/"><img src="/images/proyectos_de_gobierno/4.jpg" width="200px" target="_blank"></a>
				<!--<a href="http://distancia.ues.edu.sv/"><img src="/images/proyectos_de_gobierno/uonline.png" width="350px" target="_blank"></a>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;
		     	<a href="http://becas.rree.gob.sv/"><img src="/images/proyectos_de_gobierno/becas.jpg"  width="250px" target="_blank"></a>-->
			

			</div>
	</div>
</div>
</div>

	
			
		<main id="content" role="main" class="span6">
					<!-- Begin Content -->
					
					<div id="system-message-container">
	</div>

					
					
					<!-- End Content -->
				</main>
				
		
		</div>
		
</div> <!--FIN BODY-->
	
	<!-- Footer -->
	<footer class="footer" role="contentinfo">

		<div class="container">
<!-- 			<hr /> -->
		
							<!-- Begin Sidebar -->
					<div id="sidebar" class="span3 interes">
						<div class="sidebar-nav">
									<div class="moduletable interes">
							<h3>Lo más buscado</h3>
						<ul class="nav menu nav-pills">
<li class="item-334"><a href="/index.php/esmate" >Proyecto de Mejoramiento de Aprendizajes en Matemática en Educación Básica y Educación Media (ESMATE)</a></li><li class="item-166"><a href="/index.php/coleccion-cipotes" >Colección Cipotes</a></li><li class="item-167"><a href="http://www.mined.gob.sv/index.php/licitaciones" >Zona de Contrataciones Institucionales</a></li><li class="item-168"><a href="/index.php/directorio-centros-educativos" >Directorio Centros Educativos</a></li><li class="item-169"><a href="http://www.mined.gob.sv/index.php/descargas/category/661-colegios-privados" >Colegios privados</a></li><li class="item-170"><a href="/index.php/2015-05-12-15-21-32" >Programas de estudio</a></li><li class="item-171"><a href="/index.php/estadisticas-educativas" >Estadísticas Educativas</a></li><li class="item-172"><a href="/index.php/servicios-en-linea-mined" >Servicios en Línea MINED</a></li><li class="item-174"><a href="/index.php/2015-05-12-15-29-13" >Estadísticas Educación Superior</a></li><li class="item-254"><a href="/index.php/licitaciones" >Licitaciones</a></li><li class="item-296"><a href="/index.php/foroculturadepaz" >Foro Cultura de Paz</a></li></ul>
		</div>
	
						</div>
					</div>
					<!-- End Sidebar -->
		
							<!-- Lo mas buscado -->
					<div id="sidebar" class="span3">
						<div class="sidebar-nav">
									<div class="moduletable enlaces">
							<h3>De interés</h3>
						<ul class="nav menu nav-pills">
<li class="item-160"><a href="/index.php/titulares" >Titulares</a></li><li class="item-161"><a href="/index.php/plan-social-educativo" >Plan Social Educativo</a></li><li class="item-162"><a href="http://www.presidencia.gob.sv" >Presidencia de La República</a></li><li class="item-163"><a href="http://www.miportal.edu.sv" >Mi Portal</a></li><li class="item-164"><a href="http://programaeuro-solar.eu/" >EuroSolar</a></li><li class="item-265"><a href="/index.php/gestion-de-la-calidad" >Gestion de la Calidad</a></li><li class="item-281"><a href="/index.php/programas-sociales" >Programas  Sociales</a></li><li class="item-325"><a href="/index.php/encuesta-ciudadana" >Encuesta ciudadana</a></li><li class="item-330"><a href="/index.php/observatorio" >Observatorio Nacional del Sistema Educativo</a></li><li class="item-336"><a href="/index.php/guias-y-recursos-educacion-artistica-y-fisica" >Guías y Recursos Educación Artística y Física</a></li></ul>
		</div>
	
						</div>
					</div>
					<!-- End Buscado -->
							<div id="aside" class="span4">
				

					<!-- Begin Right Sidebar -->
							<div class="moduletable social">
							<h3>Participación Ciudadana</h3>
						<!-- BEGIN: Custom advanced (www.pluginaria.com) -->
<a name="participacion" href="http://twitter.com/MINEDelsalvador"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-twitter fa-stack-1x fa-inverse"></i>
          </span>
</a> 
<a name="participacion" href="https://www.facebook.com/MINEDelsalvador"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-facebook fa-stack-1x fa-inverse"></i>
          </span>
</a>
<a name="participacion" href="https://www.youtube.com/channel/UC7JZ4j5-dQX6j8BgaASOP_Q"/>
<span class="fa-stack fa-lg">
            <i class="fa fa-circle fa-stack-2x"></i>
            <i class="fa fa-youtube fa-stack-1x fa-inverse"></i>
          </span>
</a>

    <!-- END: Custom advanced (www.pluginaria.com) -->
		</div>
	
					<!-- End Right Sidebar -->
					<p class="copy">
						<a rel="license" href="http://creativecommons.org/licenses/by-nc-nd/4.0/"><img alt="Licencia de Creative Commons" style="border-width:0" src="https://i.creativecommons.org/l/by-nc-nd/4.0/88x31.png" /></a><br /><span xmlns:dct="http://purl.org/dc/terms/" href="http://purl.org/dc/dcmitype/InteractiveResource" property="dct:title" rel="dct:type"></span> Ministerio de Educaci&oacute;n, Gobierno de El Salvador Edificios A, Plan Maestro, Centro de Gobierno, Alameda Juan Pablo II y calle Guadalupe, San Salvador, El Salvador, Am&eacute;rica Central. Tel&eacute;fonos: +(503) 2592-2122, +(503) 2592-3117 Correo electr&oacute;nico: educacion@mined.gob.sv <p> <a style="color:white" href="/index.php/contactenos/esquema-oficinas-centrales">Mapa de Ubicaci&oacute;n</a></p></p>

					</p>
			</div>
					
	<!-- 	<div class="header-search pull-right">
			
		</div> -->
			<p class="pull-right">
					
				<!--INICIO SELLO-->
					<a rel="nofollow"  title="Estandarización de Sitios Web" href="http://estandarizacion.itiges.sv/?p=537"><center> <img alt="Estandarización de Sitios Web" width="15%" src="/images/MINED.png" ></center></a>
					
				<!--FIN SELLO-->
				<center>

				<a href="#top" style="color:#fff" id="back-top">
					
					Volver arriba				</a>
				</center>
			</p>
			
		</div>
		
	</footer>

	<script type="text/javascript">
		if (navigator.userAgent.match(/IEMobile\/10\.0/)) {
    var msViewportStyle = document.createElement("style")
 
    msViewportStyle.appendChild(
        document.createTextNode(
            "@-ms-viewport{width:auto!important}"
        )
    )
 
    document.getElementsByTagName("head")[0].appendChild(msViewportStyle)
}
	</script>
<!--Escript de Google para Estadisticas -->
<script type="text/javascript">
var gaJsHost = (("https:" == document.location.protocol) ? "https://ssl." : "http://www.");
document.write(unescape("%3Cscript src='" + gaJsHost + "google-analytics.com/ga.js' async type='text/javascript'%3E%3C/script%3E"));
</script>
<script type="text/javascript">
try {
var pageTracker = _gat._getTracker("UA-912196-1");
pageTracker._trackPageview();
} catch(err) {}</script>
<script>
</script>
</body>
</html>