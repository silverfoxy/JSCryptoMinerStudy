<!DOCTYPE html>  
<!--[if IEMobile 7 ]> <html lang="es-ES"class="no-js iem7"> <![endif]-->
<!--[if lt IE 7 ]> <html lang="es-ES" class="no-js ie6"> <![endif]-->
<!--[if IE 7 ]>    <html lang="es-ES" class="no-js ie7"> <![endif]-->
<!--[if IE 8 ]>    <html lang="es-ES" class="no-js ie8"> <![endif]-->
<!--[if (gte IE 9)|(gt IEMobile 7)|!(IEMobile)|!(IE)]><!--><html lang="es-ES" class="no-js"><!--<![endif]-->
<head>
	<meta charset="utf-8">
	<!--<meta name="viewport" content="width=device-width, initial-scale=1, user-scalable=no"/>-->
	<meta name="viewport" content="width=device-width, initial-scale=1.0, maximum-scale=1.0, minimum-scale=1.0, user-scalable=no"/>
	<meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
	
	<title>Diario El Mundo | Noticias de El Salvador y el Mundo</title>	
	<link rel="pingback" href="http://elmundo.sv/xmlrpc.php">


	
	<!-- Meta Diario El Mundo -->
		<meta name="keywords" content="Noticias, El Salvador, El Mundo, Salvador, centroamerica, America, Notas, Nota, Noticia, Periódicos, Periodicos, Arena, FMLN, Diario, el mundo el salvador, diarioelmundo">
	<meta name="description" content="Diario El Mundo - Noticias de El Salvador y el Mundo">
		
	<meta name="application-name" content="Diario El Mundo">
	<meta name="generator" content="CMS" />
	<meta name="author" content="elmundo.sv"/>
	<meta name="organization" content="Grupo Mundo">
	<meta name="application-url" content="http://www.elmundo.sv">
	<meta name="google" content="notranslate">
	<meta name="lang" content="es"></meta>
    <meta http-equiv="Content-Language" content="es" />
	<meta name="locality" content="El Salvador"></meta>
	<meta name="google-site-verification" content="_"></meta>

	<!-- Google Fonts -->
	<link href="https://fonts.googleapis.com/css?family=Adamina|Merriweather|Montserrat:100,200,300,400,500,600,700|Raleway:400,700|Roboto+Condensed:300i,400i,400,700" rel="stylesheet">


	<link rel="shorcut icon" href="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/favicon.ico">
	<script src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/js/jquery.js"></script>

		<link rel="stylesheet" href="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/js/intersticial/overlaymovil.css">
	
	<!-- wordpress head functions -->
	<link rel='dns-prefetch' href='//s.w.org' />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/elmundo.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.9.4"}};
			!function(a,b,c){function d(a,b){var c=String.fromCharCode;l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,a),0,0);var d=k.toDataURL();l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,b),0,0);var e=k.toDataURL();return d===e}function e(a){var b;if(!l||!l.fillText)return!1;switch(l.textBaseline="top",l.font="600 32px Arial",a){case"flag":return!(b=d([55356,56826,55356,56819],[55356,56826,8203,55356,56819]))&&(b=d([55356,57332,56128,56423,56128,56418,56128,56421,56128,56430,56128,56423,56128,56447],[55356,57332,8203,56128,56423,8203,56128,56418,8203,56128,56421,8203,56128,56430,8203,56128,56423,8203,56128,56447]),!b);case"emoji":return b=d([55357,56692,8205,9792,65039],[55357,56692,8203,9792,65039]),!b}return!1}function f(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var g,h,i,j,k=b.createElement("canvas"),l=k.getContext&&k.getContext("2d");for(j=Array("flag","emoji"),c.supports={everything:!0,everythingExceptFlag:!0},i=0;i<j.length;i++)c.supports[j[i]]=e(j[i]),c.supports.everything=c.supports.everything&&c.supports[j[i]],"flag"!==j[i]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[j[i]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(h=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",h,!1),a.addEventListener("load",h,!1)):(a.attachEvent("onload",h),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),g=c.source||{},g.concatemoji?f(g.concatemoji):g.wpemoji&&g.twemoji&&(f(g.twemoji),f(g.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='stylesheet' id='wp-polls-css'  href='http://elmundo.sv/wp-content/plugins/wp-polls/polls-css.css?ver=2.73.8' type='text/css' media='all' />
<style id='wp-polls-inline-css' type='text/css'>
.wp-polls .pollbar {
	margin: 1px;
	font-size: 8px;
	line-height: 10px;
	height: 10px;
	background: #24558F;
	border: 1px solid #c8c8c8;
}

</style>
<link rel='stylesheet' id='bootstrap-css'  href='http://elmundo.sv/wp-content/themes/theme_elmundosv2017/library/css/bootstrap.css?ver=1.0' type='text/css' media='all' />
<link rel='stylesheet' id='wpbs-style-css'  href='http://elmundo.sv/wp-content/themes/theme_elmundosv2017/style.css?ver=1.0' type='text/css' media='all' />
<script type='text/javascript' src='http://cdn.elmundo.sv/wp-includes/js/jquery/jquery.js?ver=1.12.4'></script>
<script type='text/javascript' src='http://cdn.elmundo.sv/wp-includes/js/jquery/jquery-migrate.min.js?ver=1.4.1'></script>
<script type='text/javascript' src='http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/library/js/bootstrap.min.js?ver=1.2'></script>
<script type='text/javascript' src='http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/library/js/scripts.js?ver=1.2'></script>
<link rel='https://api.w.org/' href='http://elmundo.sv/wp-json/' />
			<style type="text/css" media="screen">
				/**
				 * Plugin Name: Subtitles
				 * Plugin URI: http://wordpress.org/plugins/subtitles/
				 * Description: Easily add subtitles into your WordPress posts, pages, custom post types, and themes.
				 * Author: We Cobble
				 * Author URI: https://wecobble.com/
				 * Version: 2.2.0
				 * License: GNU General Public License v2 or later
				 * License URI: http://www.gnu.org/licenses/gpl-2.0.html
				 */

				/**
				 * Be explicit about this styling only applying to spans,
				 * since that's the default markup that's returned by
				 * Subtitles. If a developer overrides the default subtitles
				 * markup with another element or class, we don't want to stomp
				 * on that.
				 *
				 * @since 1.0.0
				 */
				span.entry-subtitle {
					display: block; /* Put subtitles on their own line by default. */
					font-size: 0.53333333333333em; /* Sensible scaling. It's assumed that post titles will be wrapped in heading tags. */
				}
				/**
				 * If subtitles are shown in comment areas, we'll hide them by default.
				 *
				 * @since 1.0.5
				 */
				#comments .comments-title span.entry-subtitle {
					display: none;
				}
			</style>	<!-- end of wordpress head -->

	<!-- IE8 fallback moved below head to work properly. Added respond as well. Tested to work. -->
		<!-- media-queries.js (fallback) -->
	<!--[if lt IE 9]>
		<script src="http://css3-mediaqueries-js.googlecode.com/svn/trunk/css3-mediaqueries.js"></script>			
	<![endif]-->

	<!-- html5.js -->
	<!--[if lt IE 9]>
		<script src="http://html5shim.googlecode.com/svn/trunk/html5.js"></script>
	<![endif]-->	
	
	<!-- respond.js -->
	<!--[if lt IE 9]>
          <script type='text/javascript' src="http://cdnjs.cloudflare.com/ajax/libs/respond.js/1.4.2/respond.js"></script>
	<![endif]-->

	<!-- Carrousel Clima/Boton Suscribase -->
	<link rel="stylesheet" href="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/css/jquery.bxslider.css" type="text/css" />
	<script src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/js/jquery.bxslider.js"></script>
	<script type="text/javascript">
		var j = jQuery.noConflict();
		j(document).ready(function() 
			{
			j('.bxslider').bxSlider({
			    auto: true,
				autoControls: false,
				controls: false,
				pager: false,
			    mode: 'fade',
			    pause:8000
			});
		}); 

		var fg = jQuery.noConflict();
		fg(document).ready(function() 
			{
			fg('.postslider').bxSlider({
			    auto: true,
				autoControls: false,
				controls: true,
				pager: false,
			    mode: 'fade',
			    pause:6000
			});
		});

		var vi = jQuery.noConflict();
		vi(document).ready(function() 
			{
			vi('.postslider2').bxSlider({
			    auto: true,
				autoControls: false,
				controls: true,
				pager: false,
			    mode: 'fade',
			    pause:5000
			});
		});

		//Pautas
		var pa = jQuery.noConflict();
		pa(document).ready(function() 
			{
			pa('.pautas-print').bxSlider({
			    auto: true,
				autoControls: false,
				controls: true,
				pager: false,
			    mode: 'fade',
			    pause:5000
			});
		}); 

	</script>
	<!-- Finaliza carrousel -->

<!--  ENVIVO -->
	<style>
	.box {
		display: none;
	  width: 20%;
	  margin: 0 auto;
	  background: rgba(255,255,255,0.2);
	  padding: 35px;
	  border: 2px solid #fff;
	  border-radius: 20px/50px;
	  background-clip: padding-box;
	  text-align: center;
	}

	.button {
	  font-size: 1em;
	  padding: 10px;
	  color: #fff;
	  border: 2px solid orange;
	  border-radius: 20px/50px;
	  text-decoration: none;
	  cursor: pointer;
	  transition: all 0.3s ease-out;
	}
	.button:hover {
	  background: orange;
	}


	.popup {
		padding: 5px;
		background: #444;
		border-radius: 2px;
		width: 25%;
		position: fixed;
		transition: all 0.5s ease-in-out;
		bottom: 0;
		top: auto;
		right: 0;
	}

	.popup h2 {
	  margin: 0 0 2px 0;
	  color: #fff;
	  font-size: 11px;
	  font-weight: normal;
	  font-family: Tahoma, Arial, sans-serif;
	}
	.popup .close {
	  position: absolute;
	  top: 0px;
	  right: 20px;
	  transition: all 0.5s;
	  font-size: 20px;
	  font-weight: bold;
	  text-decoration: none;
	  color: #fff;
	}
	.popup .close:hover {
	  color: red;
	}
	.popup .content {
	  max-height: 30%;
	  overflow: auto;
	}
	@media screen and (max-width: 768px) {
	    .popup {
			display: none !important;
	    }
	}
	</style>	


	<!-- Google Analytics -->
	<script>
	  (function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
	  (i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
	  m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
	  })(window,document,'script','//www.google-analytics.com/analytics.js','ga');
	
	  ga('create', 'UA-16962426-3', 'auto');
	  
	  	  //Home
	  ga('set', 'contentGroup1', 'HME');
	  	
	  	  	  	  	  	  	  	  	  	  	  	  	  	  	  
	  //*** Tracking in Google Analytics the autor post ***
	  	  //*** End traking code ***

	  ga('send', 'pageview');
	  setTimeout("ga('send','event','Permanencia','>60 segs')",60000);
	</script>


	
	<!--############################## Universal DFP #################################-->
	<script src='https://www.googletagservices.com/tag/js/gpt.js'></script>

	<script>
	  	googletag.cmd.push(function() {
	    googletag.defineSlot('/12206962/dem_sky1', [[970, 90], [320, 100]], 'div-gpt-ad-1499235990987-0').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_btn1', [220, 90], 'div-gpt-ad-1499235990987-1').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_lead1', [[320, 100], [728, 90]], 'div-gpt-ad-1499235990987-2').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_lead2', [[320, 100], [728, 90]], 'div-gpt-ad-1499235990987-3').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_rect0', [[300, 250], [600, 380]], 'div-gpt-ad-1499235990987-4').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_rect1', [300, 250], 'div-gpt-ad-1499235990987-5').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_rect2', [300, 600], 'div-gpt-ad-1499235990987-6').addService(googletag.pubads());
	    googletag.defineSlot('/12206962/dem_rect3', [[300, 600], [300, 250]], 'div-gpt-ad-1499235990987-7').addService(googletag.pubads());
	    	    		//Home
		googletag.pubads().setTargeting('dem_sec', ['HME']);
			
																														
	    googletag.pubads().enableSingleRequest();
	    googletag.pubads().collapseEmptyDivs();
	    googletag.pubads().enableSyncRendering();
	    googletag.enableServices();
	  });
	</script>
	
	<script>
		
		/*$(document).ready(function(){
			if ($('#div-gpt-ad-1498601967371-0').css('height') === '90px') {
		    	$('#div-gpt-ad-1498601967371-0').css({

		    	})
		    }else{
		    	alert('Expandir');
		    			    	Expand		    }
		});*/
		
	</script>
	<!-- Expandibles -->

	
	<style>
		
		/*------------------------------------------------------------------------------------*/
		/* Home | Publicidades | Nacionales | Economia | Entretenimiento */ 
		#div-gpt-ad-1499235990987-0{
			display: none;
		}
		#div-gpt-ad-1499235990987-0{
			background-color:#fff;
			outline: none;
			overflow: hidden!important;
			height: 90px!important;
			/* Set our transitions up. */
			-webkit-transition: all 0.8s;
			-moz-transition: all 0.8s;
			transition: all 0.8s;
		}
		#div-gpt-ad-1499235990987-0:hover{
			height: 415px!important;
		}
		#div-gpt-ad-1499235990987-0:hover iframe{
			margin-top: -90px;
		}
		
	</style>
	
	
	<!--############################## End Universal DFP #################################-->

	
	<!-- MailChimpForm -->
	<link href="http://cdn-images.mailchimp.com/embedcode/horizontal-slim-10_7.css" rel="stylesheet" type="text/css">
	<style type="text/css">
		#mc_embed_signup{background:#ececec; clear:left; width:100%;padding: 15px;margin-bottom: 20px;}

		#mc_embed_signup h3{
		    color: #555;
		    font-size: 24px;
		    letter-spacing: -1px;
		    margin: 0;
		} 
		#mc_embed_signup h3 span{
			display: block;
			color: #B90004;
		}
		#mc_embed_signup label{
			font-weight: normal;
			font-size: 12px;
			text-align: left;
		}
		#mc_embed_signup input{
			width: 100%!important;
		}
		#mc_embed_signup .clear{
			display: block!important;
			margin-top: 32px;
		}
		#mc_embed_signup .button{
			background: #B90004;
			transition:all 0.23s ease-in-out 0s;
		}
		/*#mc_embed_signup form div#mc_embed_signup_scroll div.clear input{
			width: 100%!important;
		}*/

		/* Add your own MailChimp form style overrides in your site stylesheet or in this style block.
		   We recommend moving this block and the preceding CSS link to the HEAD of your HTML file. */
	</style>
	<!-- /MailChimpForm -->

	    <!-- End Wordpres Gallery -->

	<!-- Anuncio CopaAmerica -->
	<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
	

	<link rel="stylesheet" href="https://cdnjs.cloudflare.com/ajax/libs/animate.css/3.5.2/animate.css">


	<!--script>
		var deviceDnm =  $(window).width();
		alert("Ancho: " + deviceDnm);
		
		if(deviceDnm <= 768){
			//alert("Es menor, muestro version movil");
			var wrapperMv = document.getElementById('dsDnm');
			wrapperMv.onload = function() {
			    alert("Content loaded, removing iframe...");
			    this.parentNode.removeChild(this);    
			};
			document.body.appendChild(wrapperMv);
		}else{
			//alert("Es mayor, muestro version desktop");
			var wrapperDs = document.getElementById('mvDnm');
			wrapperDs.onload = function() {
			    alert("Content loaded, removing iframe...");
			    this.parentNode.removeChild(this);    
			};
			document.body.appendChild(wrapperDs);
		}
	</script-->

	<!-- Perfect Scroll navmenu -->
	<link href="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/js/perfect-scrollbar.min.css" rel="stylesheet">

	</head>

	<body class="home blog">
		
		<!-- /12206962/dem_rect0 -->
		<div id='div-gpt-ad-1499235990987-4'>
			<div id="boxesmovil" class="">
				<div id="popupmovil" class="windowmovil">
					<div style="font-family: Arial,Helvetica,sans-serif; font-size: 14px; font-weight: bold;">  
						<a href="#" class="closepubmovil">Cerrar [X]</a>
					</div>

					<script>
					googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-4'); });
					</script>
				</div>
				<!-- Mask to cover the whole screen -->
				<div style="width: 1478px; height: 602px; display: none; opacity: 0.8;" id="maskmovil"></div>
			</div>
		</div>

		<!-- /12206962/dem_rect0 -->
		
		
		<script>
		$(document).ready(function(){
			
			/* Automatizar Expand or Not the Adserver modul */
			function showHeight( element, height ) {
			  if(height === 90 || height === 100){
			  	$( "#medidaExp" ).text( "No Expand, the div is " + height + "px." );
			  	//$(this).prev('#div-gpt-ad-1498601967371-0').prop('id', 'div-gpt-ad-1498601967371-777');	
			  	$("#div-gpt-ad-1499235990987-0").prop('id', 'div-gpt-ad-1499235990987-777');
			  }else{
			  	$( "#medidaExp" ).text( "Expand, the div is " + height + "px." );
			  	$("#div-gpt-ad-1499235990987-777").prop('id', 'div-gpt-ad-1499235990987-0');
			  }
			}
			jQuery(window).on("load", function(){
				showHeight( "document", $( "#div-gpt-ad-1499235990987-0_ad_container > ins" ).height() );
				$("#div-gpt-ad-1499235990987-0").show();
			});
			/* /Automatizar Expand or Not the Adserver modul */


		    //Universal Overlay
		    if ($('#div-gpt-ad-1499235990987-4').css('display') !== 'none') {
		    	//alert('Tengo anuncio');
		    	//Inicializamos condicion movil
                /*$(document).ready(function() {
                        loadpopmovil();
                });*/
				
				setTimeout(function() { 
					loadpopmovil();
				}, 5000);

                //Funcion para mostrar Publicidad
                function loadpopmovil(){
                  var idmovil = '#popupmovil';

                  //Get the screen height and width
                  var maskHeightm = $(document).height();
                  var maskWidthm = $(window).width();

                  //Set heigth and width to mask to fill up the whole screen
                  $('#maskmovil').css({'width':maskWidthm,'height':maskHeightm});

                  //transition effect
                  $('#maskmovil').fadeIn(1000);
                  $('#maskmovil').fadeTo("slow",0.8);

                  //Get the window height and width
                  var winHm = $(window).height();
                  var winWm = $(window).width();

                  //Set the popupmovil window to center
                  $(idmovil).css('top',  winHm/2-$(idmovil).height()/2);
                  $(idmovil).css('left', winWm/2-$(idmovil).width()/2);

                  //transition effect
                  $(idmovil).fadeIn(2000);

                  setTimeout(function() { 
                    $(".closepubmovil").trigger("click");
                  }, 5000);

                  //if close button is clicked
                  $('.closepubmovil').click(function (e) {
                    //Cancel the link behavior
                    e.preventDefault();

                    $('#maskmovil').hide();
                    $('.windowmovil').hide();
                  });

                }
		    } //Cerramos el if display:none

		});
		</script>
		




		
		<!-- Menu Movil -->
		<nav class="navbar navbar-fixed-top hidden-md hidden-lg">
				
				<div class="container-fluid container-tablet-menu">
			    <!-- Brand and toggle get grouped for better mobile display -->
			    <div class="navbar-header navbar-movil2 header-tablet-menu" style="padding-bottom:5px; min-height:45px; border-bottom:2px solid #fff;">
			      <!-- Logo Movil -->
			      <!--iframe src="http://dinamo.click/index.php?l=100003" style="width:234px; height:30px; float:left!important;" width="100%" height="30" scrolling="no" frameborder="0" target="_top"></iframe-->
				  <a class="navbar-brand" href="http://elmundo.sv" style="float:left!important; margin-top:-2px;">
			      	<img src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/images/brand-dem-movil.png" alt="" class="img-responsive">
			      </a>
			      
			      <!--button type="button" class="navbar-toggle collapsed btn-menumovil" data-toggle="collapse" data-target="#bs-example-navbar-collapse-1" aria-expanded="false" style="margin-right:0; margin-top:6px; background:transparent!important;">
			        <div style="float:right;">
				        <span class="sr-only">Toggle navigation</span>
				        <span class="icon-bar"></span>
				        <span class="icon-bar"></span>
				        <span class="icon-bar"></span>
					</div>
					<div style="float:left; margin-right:12px; font-size:13px; font-weight:bold; display:none;">
			        	<span>MENÚ</span>
			        </div>
			        <div style="clear:both; overflow:hidden;"></div>
			      </button-->

			      <div class="spinner-master navbar-toggle collapsed btn-menumovil" data-toggle="collapse" data-target="#bs-example-navbar-collapse-1" aria-expanded="false" style="margin-right:0; margin-top:6px; background:transparent!important;">
					  <input type="checkbox" id="spinner-form" />
					  <label for="spinner-form" class="spinner-spin">
					    <div class="spinner diagonal part-1"></div>
					    <div class="spinner horizontal"></div>
					    <div class="spinner diagonal part-2"></div>
					  </label>
					</div>

			    </div>

			    <!-- Collect the nav links, forms, and other content for toggling -->
			    <div class="collapse navbar-collapse items-menumovil collapse-tablet-menu" id="bs-example-navbar-collapse-1" style="padding:0!important;">
  					<div class="menu-menu-principal-sin-submenu-container"><ul id="menu-menu-principal-sin-submenu" class="menu"><li id="menu-item-798364" class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-798364 active"><a href="http://elmundo.sv/">Inicio</a></li>
<li id="menu-item-632441" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632441"><a href="http://elmundo.sv/category/confidencial-editorial/">Confidencial &#038; Editorial</a></li>
<li id="menu-item-632442" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632442"><a href="http://elmundo.sv/category/nacionales/">Nacionales</a></li>
<li id="menu-item-632444" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632444"><a href="http://elmundo.sv/category/deportes/">Deportes</a></li>
<li id="menu-item-632445" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632445"><a href="http://elmundo.sv/category/entretenimiento/">Entretenimiento</a></li>
<li id="menu-item-632443" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632443"><a href="http://elmundo.sv/category/politica/">Política</a></li>
<li id="menu-item-632449" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632449"><a href="http://elmundo.sv/category/internacionales/">Internacionales</a></li>
<li id="menu-item-645514" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-645514"><a href="http://elmundo.sv/category/conectados/">Conectados</a></li>
<li id="menu-item-793738" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793738"><a href="http://elmundo.sv/category/mujer-salud/">Mujer &amp; Salud</a></li>
<li id="menu-item-632448" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632448"><a href="http://elmundo.sv/category/economia/">Economía</a></li>
<li id="menu-item-793737" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793737"><a href="http://elmundo.sv/category/empresarial/">Empresarial</a></li>
<li id="menu-item-632493" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632493"><a href="http://elmundo.sv/category/perfiles-bloggers/">Blog</a></li>
</ul></div>  					<div class="col-xs-12 buscardormovil" style="padding-bottom:8px; display:none;">
  					  					</div>
					<div class="sharedNetsMovil">
						<a href="https://www.facebook.com/ElMundoSV" target="_blank">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-facebook.svg" alt=""></a>
						<a href="http://twitter.com/ElMundoSV" target="_blank">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-twitter.svg" alt=""></a>
						<a href="https://www.linkedin.com/company/elmundosv" target="_blank">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-linkedin.svg" alt=""></a>
						<a href="https://www.youtube.com/user/DiarioElMundoTV" target="_blank">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-youtube.svg" alt=""></a>
						<a href="http://instagram.com/ElMundoSV" target="_blank">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-instagram.svg" alt=""></a>
						<a  href="http://elmundo.sv/newsletter/">
							<img width="32" height="32" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-mailw.svg" alt=""></a>
					</div>
  					<div class="col-xs-12 botonera-movil" style="text-align:right; padding-top:6px; padding-bottom:7px; border-top:1px solid rgba(36,46,56,0.85);;">
																			<a href="https://issuu.com/elmundocomsv/docs/mundo190318" target="_blank">
								E-paper <img src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/images/btn-nepaper.png" alt="">
							</a>
						
						<!--a href="http://elmundo.sv/newsletter/">
							Suscribase <img src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/images/btn-nemail.png" alt="">
						</a-->

  					</div>
				</div><!-- /.navbar-collapse -->
		  	</div><!-- /.container-fluid -->
		</nav>
		<div id="mobile-nav-wrapper" class="hidden" style="display:none;">
						</div>
		<!-- /End Menu -->

		
		<div class="container">
			<!-- LEADERBOARD -->
			
		<div id="stickyBar" >
			<!-- Logo / Main Menú -->
			<div class="row"  style='display:block;'>
				<div class="col-sm-12" style="text-align:center; padding-top:15px;">
					
					<!--
					50 Años Diario El Mundo
					position:relative; min-height:52px; DIV
					position:absolute; IMG 438 width
					-->
					<div class="hidden-xs hidden-sm visible-md visible-lg logo-tablet" style="position:relative; min-height:52px;">
					<iframe src="http://dinamo.click/index.php?l=100004" style="width:100%; height:37px" width="100%" height="37" scrolling="no" frameborder="0" target="_top"></iframe>
					</div>
					

					<a style="display:none;" href="http://elmundo.sv" class=""><img src="http://cdn.elmundo.sv/wp-content/themes/wp_bs/images/logo.png" width="438" height="51" class="img-responsive" alt="Diario El Mundo Home" title="Diario El Mundo | Sitio web de noticias e informacion para El Salvador"></a>

					<p class="date" style="margin-top:-14px;">
						
						<span style="font-weight:normal; font-size:11px;text-transform:uppercase">
							<script type="text/javascript"><!--
			                    dows = new Array("Domingo","Lunes","Martes","Mi&eacute;rcoles","Jueves","Viernes","S&aacute;bado");
			                    months = new Array("Enero","Febrero","Marzo","Abril","Mayo","Junio","Julio","Agosto","Septiembre","Octubre","Noviembre","Diciembre");

			                    now = new Date();
			                    dow = now.getDay();
			                    d = now.getDate();
			                    m = now.getMonth();
			                    h = now.getTime();
			                    y = now.getFullYear();

			                    document.write(dows[dow]+" "+d+" de "+months[m]+" de "+ y);

		                    //--></script>
						</span>
					</p>
				</div>
			</div>
			
			<div class="row"  style='display:block;'>
				<!-- Products elmundo.sv -->
				<div class="col-xs-12">
					<div class="hidden-xs hidden-sm visible-md visible-lg text-center" style="margin-bottom: 1px; margin-top:4px;">
						<div class="menu-menu-secundario-container"><ul id="menu-menu-secundario" class="menu_secundario"><li id="menu-item-701314" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-701314"><a href="http://elmundo.sv/newsletter/">Newsletter</a></li>
<li id="menu-item-793600" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-793600"><a href="http://elmundo.sv/kiosko-digital/">Kiosko Digital</a></li>
<li id="menu-item-632437" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-632437"><a href="http://vidasana.sv">VidaSana</a></li>
<li id="menu-item-632438" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-632438"><a href="http://devacaciones.sv">DeVacaciones</a></li>
<li id="menu-item-632439" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-632439"><a href="http://sanmiguel.sv/">El Migueleño</a></li>
<li id="menu-item-632440" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-632440"><a href="/especiales-diario-el-mundo/">Especiales</a></li>
<li id="menu-item-824999" class="menu-item menu-item-type-custom menu-item-object-custom menu-item-824999"><a target="_blank" href="http://mimundo.sv">Mundo Universitario</a></li>
</ul></div>					</div>
				</div>
			</div>

			<div class="row">
				<div class="col-xs-12">
					<nav class="navbar navbar-default hidden-xs hidden-sm" role="navigation" id="menu_principal" style="margin-bottom:0; border-bottom:1px solid #f4f4f4 !important">
					    <button class="hamburger">
					    	<div class="HmbBtn">
					    	<span class="linesHmb"></span>
					    	<span class="linesHmb"></span>
					    	<span class="linesHmb"></span>
					    	</div>
					    </button>
  						<button class="cross">
							<div class="CloseBtn">
  								<span>x</span>
  							</div>
  						</button>
  						<!-- BUTTONS -->
  						<!--a href="http://elmundo.sv" class="btnHomepage">INICIO</a-->
  						<!-- Button trigger searchForm -->
						<button type="button" class="btn btn-primary btnSearch" data-toggle="modal" data-target=".bs-example-modal-sm">
						</button>
						<!-- /BUTTONS -->
						

  						<div id="wrapMenu"><div class="menu-menu-principal-sin-submenu-container"><ul id="menu-menu-principal-sin-submenu-1" class="hamburgerMenu perfectScroll"><li class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-798364 active"><a href="http://elmundo.sv/">Inicio</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632441"><a href="http://elmundo.sv/category/confidencial-editorial/">Confidencial &#038; Editorial</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632442"><a href="http://elmundo.sv/category/nacionales/">Nacionales</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632444"><a href="http://elmundo.sv/category/deportes/">Deportes</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632445"><a href="http://elmundo.sv/category/entretenimiento/">Entretenimiento</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632443"><a href="http://elmundo.sv/category/politica/">Política</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632449"><a href="http://elmundo.sv/category/internacionales/">Internacionales</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-645514"><a href="http://elmundo.sv/category/conectados/">Conectados</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793738"><a href="http://elmundo.sv/category/mujer-salud/">Mujer &amp; Salud</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632448"><a href="http://elmundo.sv/category/economia/">Economía</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793737"><a href="http://elmundo.sv/category/empresarial/">Empresarial</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632493"><a href="http://elmundo.sv/category/perfiles-bloggers/">Blog</a></li>
</ul></div>						<div class="sharedNets">
							<a href="https://www.facebook.com/ElMundoSV" target="_blank">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-facebook.svg" alt=""></a>
							<a href="http://twitter.com/ElMundoSV" target="_blank">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-twitter.svg" alt=""></a>
							<a href="https://www.linkedin.com/company/elmundosv" target="_blank">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-linkedin.svg" alt=""></a>
							<a href="https://www.youtube.com/user/DiarioElMundoTV" target="_blank">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-youtube.svg" alt=""></a>
							<a href="http://instagram.com/ElMundoSV" target="_blank">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-instagram.svg" alt=""></a>
							<a href="http://elmundo.sv/newsletter/">
								<img width="28" height="28" src="http://elmundo.sv/wp-content/themes/theme_elmundosv2017/images/ico-mail.svg" alt=""></a>
						</div>
						</div>

					    <div id="wrapNav" class="container-fluid">

				    		<div id="nav_menu-2" class="widget widget_nav_menu main-menu"><div class="menu-menu-principal-sin-submenu-container"><ul id="menu-menu-principal-sin-submenu-2" class="menu"><li class="menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home menu-item-798364 active"><a href="http://elmundo.sv/">Inicio</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632441"><a href="http://elmundo.sv/category/confidencial-editorial/">Confidencial &#038; Editorial</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632442"><a href="http://elmundo.sv/category/nacionales/">Nacionales</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632444"><a href="http://elmundo.sv/category/deportes/">Deportes</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632445"><a href="http://elmundo.sv/category/entretenimiento/">Entretenimiento</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632443"><a href="http://elmundo.sv/category/politica/">Política</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632449"><a href="http://elmundo.sv/category/internacionales/">Internacionales</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-645514"><a href="http://elmundo.sv/category/conectados/">Conectados</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793738"><a href="http://elmundo.sv/category/mujer-salud/">Mujer &amp; Salud</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632448"><a href="http://elmundo.sv/category/economia/">Economía</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-793737"><a href="http://elmundo.sv/category/empresarial/">Empresarial</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-632493"><a href="http://elmundo.sv/category/perfiles-bloggers/">Blog</a></li>
</ul></div></div>

					    </div><!-- /.container-fluid -->
						<div id="imgBrand">
					    	<a href="http://elmundo.sv">
					    		<img src="http://static.elmundo.sv/wp-content/uploads/2017/10/dem-lred.png" alt="">
					    	</a>
					    </div>
					    <!--div id="searchBrand">
					    						    </div-->
					</nav>
				</div>

			</div>

		</div>


		<!-- ========= Skyscraper Ad =============== -->
					<div class="row" style="text-align:center;">
				<div class="col-xs-12 moveTopDsk">
					<div class="adblockweb" style="text-align:center;">
	<div id="text-52" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_sky1 -->
<div id='div-gpt-ad-1499235990987-0'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-0'); });
</script>
</div></div>
		</div></div>					<script type="text/javascript">

						$(document).ready(function () {

							$('#div-gpt-ad-1498160898700-4').hover(
								function () {
									$(this).stop(true, false).animate({ opacity: 1.0, width:970+'px', height: 402+'px'}, 550)
								}, 
								function () {
									$(this).stop(true, false).animate({ opacity: 1.0, width:970+'px', height:  90+'px'}, 550)
								}
							);
						});
					</script>
				</div>
			</div>
		
</div>

			
			

<script type="text/javascript">
	$(document).ready(function(){
		$("#wunderground_forecast_widget-2 .wu-copyright").hide();
		$("#wunderground_forecast_widget-2 .wu-cond-low").hide();
		$(".wu-wrapper table *").css("font-size","10px");
		$("#wunderground_forecast_widget-2 .wu-wrapper").css({'height':'90px','margin-top':'-20px'});
		$("#wunderground_forecast_widget-2").css('padding-left','18px').css('background','#134A73');
		$("#wunderground_forecast_widget-2 .wu-wrapper .wu-icon").css("margin-bottom",'0');
		$("#wunderground_forecast_widget-2 .wu-wrapper .wu-icon img").css({'height':'40px','width':'40px'});
		$("#wunderground_forecast_widget-2 .wu-forecast-wrapper .wu-cond-highlow").css('margin-top','2px').css('white-space','nowrap');
		$("#wunderground_forecast_widget-2 .wu-forecast-header").css("margin",'0px');
		$("#wunderground_forecast_widget-2 .wu-table-3 thead").hide();
	});
</script>

<div class="container">

	<!-- Nota en Desarrollo -->
    <div class="row">
    	<div id="execphp-10" class="widget widget_execphp">			<div class="execphpwidget"><br>
</div>
		</div>    </div>

	<div class="separator"></div>

	<div class="row" style="margin-left:0!important; margin-right:0!important;">
		<div class="col-xs-12 col-sm-12 col-md-9 col-lg-9 nopadding BreakingNews">
			<!-- RECENT POST FROM ALL CATEGORIES -->
					
									<!-- Inicia Row -->
			<div class="row">
		        <div class="col-xs-12 col-sm-8 col-md-8">
		        	<h1 class="mainHeaders moveTitle"><span>Actualidad</span></h1>
					<div class="main-thumbnail">
						<!-- Imagen destacada o primer imagen del post -->
						<a href="http://elmundo.sv/equipo-de-fuera-de-juego-vencio-al-magico-y-sus-amigos/" class="thumbnail-wrapper">
						<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Fuera-de-Juego1.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
							<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Fuera-de-Juego1.jpg" class="img-responsive thumbnail-wrapper" style="width:100%;"-->
												</a>

					</div>
		        
			        <div class="col-xs-12 nopadding">
						<h1 class="MainTitleHeader"><a href="http://elmundo.sv/equipo-de-fuera-de-juego-vencio-al-magico-y-sus-amigos/">Equipo de Fuera de Juego venció al “Mágico” y sus amigos</a></h1>
						<p>

El combinado del programa Fuera de Juego de ESPN derrotó esta tarde en la vía …</p>					</div>
				</div>
			
							<div class="col-xs-12 col-sm-4 col-md-4">
					<div class="main-thumbnail">
						
						<!-- Imagen destacada o primer imagen del post -->
						<a href="http://elmundo.sv/mourinho-pone-40-millones-por-un-consentido-de-zidane/" class="thumbnail-wrapper">
						<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Mourinho-Florentino.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
						<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Mourinho-Florentino.jpg" class="img-responsive thumbnail-wrapper"-->
												</a>

					</div>
					<h1 class="SecondTitleHeader"><a href="http://elmundo.sv/mourinho-pone-40-millones-por-un-consentido-de-zidane/">Mourinho pone $40 millones por un consentido de Zidane</a></h1>
				</div>
							<div class="col-xs-12 col-sm-4 col-md-4">
					<div class="main-thumbnail">
						
						<!-- Imagen destacada o primer imagen del post -->
						<a href="http://elmundo.sv/pupusas-de-olocuilta-obtienen-proteccion-de-propiedad-intelectual/" class="thumbnail-wrapper">
						<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Pupusas2.png" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
						<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Pupusas.png" class="img-responsive thumbnail-wrapper"-->
												</a>

					</div>
					<h1 class="SecondTitleHeader"><a href="http://elmundo.sv/pupusas-de-olocuilta-obtienen-proteccion-de-propiedad-intelectual/">Pupusas de Olocuilta obtienen protección de propiedad intelectual</a></h1>
				</div>
			<!-- Finaliza Row -->
			</div>
						<!-- Inicia Row nuevamente -->
			<div class="row">
				<div class="col-xs-12 col-sm-4 col-md-4">
					<div class="main-thumbnail">
						<!-- Imagen destacada o primer imagen del post -->
						<a href="http://elmundo.sv/fbi-infiltro-a-la-ms-13-en-estados-unidos/" class="thumbnail-wrapper">
						<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/MS-13.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
						<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/MS-13.jpg" class="img-responsive thumbnail-wrapper"-->
												</a>

					</div>
					<h1 class="SecondTitleHeader"><a href="http://elmundo.sv/fbi-infiltro-a-la-ms-13-en-estados-unidos/">FBI infiltró a la MS-13 en Estados Unidos</a></h1>
					<p>

El Buró Federal de Investigaciones (FBI) ha logrado convencer a miembros de la Mara Salvatrucha (MS-13) …</p>				</div>
							<div class="col-xs-12 col-sm-4 col-md-4">
					<div class="main-thumbnail">
						<!-- Imagen destacada o primer imagen del post -->
						<a href="http://elmundo.sv/medico-denuncia-que-en-hospital-zacamil-no-hay-ni-jeringas/" class="thumbnail-wrapper">
						<img src="http://static.elmundo.sv/wp-content/uploads/2018/01/Hospital-Zacamil.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
						<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/01/Hospital-Zacamil.jpg" class="img-responsive thumbnail-wrapper"-->
												</a>

					</div>
					<h1 class="SecondTitleHeader"><a href="http://elmundo.sv/medico-denuncia-que-en-hospital-zacamil-no-hay-ni-jeringas/">Médico denuncia que en hospital Zacamil no hay ni jeringas</a></h1>
					<p>
El médico, Carlos Ramos Hinds, reveló las carencias por las que pasa el hospital Zacamil, en …</p>				</div>
							<div class="col-xs-12 col-sm-4 col-md-4">
					<div class="SpecialBox">
						<h1 class="HeaderEnterese"><span>ENTÉRESE</span></h1>
						<div class="col-xs-12 nopadding">
							<div class="col-xs-4 nopadding">
								<div class="main-thumbnail">
									<!-- Imagen destacada o primer imagen del post -->
									<a href="http://elmundo.sv/mister-chip-al-alianza-justo-hasta-ahi-llego-el-real-madrid-de-zidane/" class="thumbnail-wrapper">
									<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/alianza2.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
									<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/alianza2.jpg" class="img-responsive thumbnail-wrapper"-->
																		</a>
								</div>
							</div>
							<div class="col-xs-8">				
								<h1 class="ThirdTitleHeader"><a href="http://elmundo.sv/mister-chip-al-alianza-justo-hasta-ahi-llego-el-real-madrid-de-zidane/">Míster Chip al Alianza: “Justo hasta ahí llegó el Real Madrid de Zidane”</a></h1>
							</div>
						</div>
				<span class="separatorPost"></span>
							<div class="col-xs-12 nopadding">
					<div class="col-xs-4 nopadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/ee-uu-sanciona-a-otros-cuatro-venezolanos-vinculados-al-gobierno/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/TRUMP3.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
							<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/TRUMP3.jpg" class="img-responsive thumbnail-wrapper"-->
														</a>
						</div>
					</div>
					<div class="col-xs-8">				
						<h1 class="ThirdTitleHeader"><a href="http://elmundo.sv/ee-uu-sanciona-a-otros-cuatro-venezolanos-vinculados-al-gobierno/">EE.UU. sanciona a otros cuatro venezolanos vinculados al gobierno</a></h1>
					</div>
				</div>
				<span class="separatorPost"></span>
							<div class="col-xs-12 nopadding">
					<div class="col-xs-4 nopadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/presidente-anuncia-cambios-en-hacienda-minec-anda-y-migracion/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/presidente.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
							<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/presidente.jpg" class="img-responsive thumbnail-wrapper"-->
														</a>

						</div>
					</div>
					<div class="col-xs-8">				
						<h1 class="ThirdTitleHeader"><a href="http://elmundo.sv/presidente-anuncia-cambios-en-hacienda-minec-anda-y-migracion/">Presidente hace ocho cambios en su gabinete</a></h1>
					</div>
					<div class="separador"></div>
				</div>
				<div class="clear"></div>
			</div>
			</div>
			<div class="col-xs-12 visible-xs visible-sm visible-md hidden-lg"><hr class="clear"></div>
			</div>
												<!-- /RECENT POST FROM ALL CATEGORIES -->
			
		</div>
		<div class="col-xs-12 col-sm-12 col-md-3 col-lg-3">
			<div class="col-xs-12 nopadding widget" id="MundoDigital">
				<!--h3 class="widgettitle">El Mundo TV</h3-->
				<div class="video-container" style="width: 100%; min-height:165px">
				<iframe src="https://www.youtube.com/embed/WlW3bH5XHCc" frameborder="0" allowfullscreen></iframe>
			  <div class="clear"></div></div><br /><div id="text-60" class="widget widget_text">			<div class="textwidget"><div id="multimedia-dem">
<h3>Suscr&iacute;base a nuestro canal</h3>
</div>
<script src="https://apis.google.com/js/platform.js"></script>
<div class="g-ytsubscribe" data-channel="DiarioElMundoTV" data-layout="full" data-count="undefined"></div></div>
		</div>			</div>
			
			<div class="col-xs-12 col-sm-6 col-md-12 nopadding widget">
				<div class="adblockweb" style="text-align:center;">
	<div id="text-57" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_rect1 -->
<div id='div-gpt-ad-1499235990987-5' style='height:250px; width:300px;'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-5'); });
</script>
</div></div>
		</div></div>			</div>
			
			<div class="col-xs-12 col-sm-6 col-md-12 widget moreRead">
				<div id="mostreadpostswidget-6" class="widget widget_mostreadpostswidget"><h2 class="widgettitle">Top 5 | Lo más leído</h2>
<table class="mlrp_ul"><tr><td><span class="top5_number">1</span></td><td><a title="Sánchez Cerén anunciaría hoy cambios en gabinete" href="http://elmundo.sv/sanchez-ceren-anunciaria-hoy-cambios-en-gabinete/"><img width="128" height="73" src="http://static.elmundo.sv/wp-content/uploads/2018/03/Consejo-de-ministros.jpg" class="attachment-thumbnail size-thumbnail" alt="" /></a></td><td><a title="Sánchez Cerén anunciaría hoy cambios en gabinete" href="http://elmundo.sv/sanchez-ceren-anunciaria-hoy-cambios-en-gabinete/"><p><span class="category_name">Sánchez Cerén anunciaría hoy cambios en gabinete</span></p></a><p style="display:none;"></p></td></tr><tr><td><span class="top5_number">2</span></td><td><a title="Presidente hace ocho cambios en su gabinete" href="http://elmundo.sv/presidente-anuncia-cambios-en-hacienda-minec-anda-y-migracion/"><img width="128" height="73" src="http://static.elmundo.sv/wp-content/uploads/2018/03/presidente.jpg" class="attachment-thumbnail size-thumbnail" alt="" /></a></td><td><a title="Presidente hace ocho cambios en su gabinete" href="http://elmundo.sv/presidente-anuncia-cambios-en-hacienda-minec-anda-y-migracion/"><p><span class="category_name">Presidente hace ocho cambios en su gabinete</span></p></a><p style="display:none;"></p></td></tr><tr><td><span class="top5_number">3</span></td><td><a title="Así reaccionó Eugenio Chicas tras ser removido del gabinete de Gobierno" href="http://elmundo.sv/asi-reacciono-eugenio-chicas-tras-ser-removido-del-gabinete-de-gobierno/"><img width="128" height="73" src="http://static.elmundo.sv/wp-content/uploads/2017/05/Eugenio-Chicas2.jpg" class="attachment-thumbnail size-thumbnail" alt="" /></a></td><td><a title="Así reaccionó Eugenio Chicas tras ser removido del gabinete de Gobierno" href="http://elmundo.sv/asi-reacciono-eugenio-chicas-tras-ser-removido-del-gabinete-de-gobierno/"><p><span class="category_name">Así reaccionó Eugenio Chicas tras ser removido del gabinete de Gobierno</span></p></a><p style="display:none;"></p></td></tr><tr><td><span class="top5_number">4</span></td><td><a title="Presentadores de ESPN y Amigos del Mágico jugarán en el ‘Cusca’" href="http://elmundo.sv/presentadores-de-espn-y-amigos-del-magico-jugaran-en-el-cusca/"><img width="128" height="73" src="http://static.elmundo.sv/wp-content/uploads/2018/03/Magico-Gonzalez-2.jpg" class="attachment-thumbnail size-thumbnail" alt="" /></a></td><td><a title="Presentadores de ESPN y Amigos del Mágico jugarán en el ‘Cusca’" href="http://elmundo.sv/presentadores-de-espn-y-amigos-del-magico-jugaran-en-el-cusca/"><p><span class="category_name">Presentadores de ESPN y Amigos del Mágico jugarán en el ‘Cusca’</span></p></a><p style="display:none;"></p></td></tr><tr><td><span class="top5_number">5</span></td><td><a title="“Lo que no se tolera al FMLN es la actitud con la corrupción”" href="http://elmundo.sv/lo-que-no-se-tolera-al-fmln-es-la-actitud-con-la-corrupcion/"><img width="128" height="73" src="http://static.elmundo.sv/wp-content/uploads/2018/03/Salvador-Samayoa.jpg" class="attachment-thumbnail size-thumbnail" alt="" /></a></td><td><a title="“Lo que no se tolera al FMLN es la actitud con la corrupción”" href="http://elmundo.sv/lo-que-no-se-tolera-al-fmln-es-la-actitud-con-la-corrupcion/"><p><span class="category_name">“Lo que no se tolera al FMLN es la actitud con la corrupción”</span></p></a><p style="display:none;"></p></td></tr></table>
		<div style="clear:both;"></div></div>			</div>
			
		</div>
	</div>
	
	<div class="clear separador"></div>
	
	<div class="row">
		<!-- Leaderboard  -->
		<div class="col-xs-12 col-sm-12 col-md-9 text-center" style="">
			<div class="ad">
			 <div class="adblockweb" style="text-align:center;">
	<div id="text-54" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_lead1 -->
<div id='div-gpt-ad-1499235990987-2'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-2'); });
</script>
</div></div>
		</div></div>	
			</div>
		</div>
		<div class="col-xs-12 col-sm-12 col-md-3 text-center" style="">
			<div class="ad">
			 <div class="adblockweb" style="text-align:center;">
	<div id="text-53" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_btn1 -->
<div id='div-gpt-ad-1499235990987-1' style='height:90px; width:220px; margin:0 auto;'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-1'); });
</script>
</div></div>
		</div><div id="execphp-14" class="widget widget_execphp">			<div class="execphpwidget"></div>
		</div></div>	
			</div>
		</div>
	</div>

	<div class="clear sepadador"></div>


	<div class="row" style="margin-left:0!important; margin-right:0!important;">
		<!-- Post Category Column -->
		<div class="col-xs-12 col-sm-12 col-md-9 nopadding">
			<!-- Videos -->
			<!--iframe 
	width="100%" 
	frameborder="0" 
	scrolling="no" 
	src="http://elmundo.sv/mundomediapp/index.php" 
	onload="this.style.height=this.contentDocument.body.scrollHeight +'px';">
</iframe-->
<iframe width="100%" frameborder="0" 
	scrolling="no" 
	id="result" 
	height="264" 
	src="http://elmundo.sv/mundomediapp/index.php">
</iframe>			<!--/Videos -->			
			
			<div class="clear"></div>
			<!--/Videos -->

			<div class="separador"></div>

			<!-- Block Post -->
			<div class="col-xs-12 nopadding boxCategories">
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/nacionales">
							NACIONALES
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/un-herido-deja-ataque-armado-en-calle-concepcion/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/taller.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/taller.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/un-herido-deja-ataque-armado-en-calle-concepcion/">Un herido deja ataque armado en Calle Concepción</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/a-estos-medicos-el-minsal-debe-el-pago-de-tres-meses/">A estos médicos el Minsal debe el pago de tres meses</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/mas-de-diez-personas-perdieron-la-vida-este-fin-de-semana-en-accidentes-de-transito/">Más de diez personas perdieron la vida este fin de semana en accidentes de tránsito </a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<div class="dotsBottom"></div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/deportes">
							DEPORTES
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/antonella-publica-tierna-fotografia-de-messi-con-sus-3-hijos-por-dia-del-padre/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/messi2.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/messi2.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/antonella-publica-tierna-fotografia-de-messi-con-sus-3-hijos-por-dia-del-padre/">Antonella publica tierna fotografía de Messi con sus 3 hijos por Día del Padre</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/presentadores-de-espn-y-amigos-del-magico-jugaran-en-el-cusca/">Presentadores de ESPN y Amigos del Mágico jugarán en el ‘Cusca’</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/rakitic-avisa-la-salida-de-un-intocable-de-florentino-perez-y-sus-cinco-pretendientes/">Rakitic avisa la salida de un “intocable” de Florentino Pérez y sus cinco pretendientes</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<div class="dotsBottom"></div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/entretenimiento">
								ENTRETENIMIENTO
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/asi-comienza-el-verano-la-ex-miss-mundo-el-salvador/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/miss-2.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/miss-2.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/asi-comienza-el-verano-la-ex-miss-mundo-el-salvador/">Así comienza el verano la ex Miss Mundo El Salvador</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/blac-chyna-envio-un-mensaje-a-rob-kardashian-por-su-cumpleanos/">Blac Chyna envío un mensaje a Rob Kardashian por su cumpleaños</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/esta-es-la-reaccion-de-angelina-jolie-al-ver-que-esta-envejeciendo/">Esta es la reacción de Angelina Jolie al ver que está envejeciendo</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/politica">
								POLÍTICA
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/asi-reacciono-eugenio-chicas-tras-ser-removido-del-gabinete-de-gobierno/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2017/05/Eugenio-Chicas2.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2017/05/Eugenio-Chicas2.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/asi-reacciono-eugenio-chicas-tras-ser-removido-del-gabinete-de-gobierno/">Así reaccionó Eugenio Chicas tras ser removido del gabinete de Gobierno</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/polemica-por-representantes-de-coalicion-arena-pcn-retrasa-conteo-de-san-vicente/">Polémica por representantes de coalición ARENA-PCN retrasa conteo de San Vicente</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/asi-quedaran-las-posiciones-en-papeleta-para-elegir-candidato-presidencial-de-arena/">Así quedarán las posiciones en papeleta para elegir candidato presidencial de ARENA</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/internacionales">
								INTERNACIONAL
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/nicaraguenses-protestan-ante-intento-de-gobierno-de-controlar-redes-sociales/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Nicaragua-Redes-Sociales.png" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Nicaragua-Redes-Sociales.png" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/nicaraguenses-protestan-ante-intento-de-gobierno-de-controlar-redes-sociales/">Nicaragüenses protestan ante intento de gobierno de controlar redes sociales</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/al-menos-un-herido-por-balacera-en-turistica-plaza-comercial-de-mexico/">Al menos un herido por balacera en turística plaza comercial de México</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/guatemala-extiende-por-seis-meses-alerta-por-sarampion/">Guatemala extiende por seis meses alerta por sarampión</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/conectados">
								CONECTADOS
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/facebook-sacudido-por-escandalo-de-violacion-de-datos-personales/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2017/11/moderadorfacebook.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2017/11/moderadorfacebook.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/facebook-sacudido-por-escandalo-de-violacion-de-datos-personales/">Facebook sacudido por escándalo de violación de datos personales</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/el-cambio-climatico-causara-una-catastrofe-migratoria-advierte-el-banco-mundial/">El cambio climático causará una catástrofe migratoria, advierte el Banco Mundial</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/madres-cantan-junto-a-sus-hijos-con-sindrome-de-down-en-emotivo-video/">Madres cantan junto a sus hijos con síndrome de Down en emotivo video</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/mujer-salud">
								MUJER & SALUD
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/esta-enfermedad-es-la-segunda-causa-de-ceguera-en-el-mundo/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/ojos1.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/ojos1.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/esta-enfermedad-es-la-segunda-causa-de-ceguera-en-el-mundo/">Esta enfermedad es la segunda causa de ceguera en el mundo</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/lo-que-no-debes-decir-a-tu-pareja-sobre-tus-ex/">Lo que no debes decir a tu pareja sobre tus ex</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/fiebre-tifoidea-como-evitarla/">Fiebre Tifoidea: ¿Cómo evitarla?</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/economia">
								ECONOMÍA
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/plaza-marinera-estaria-lista-en-primer-trimestre-de-2019/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2017/09/Puerto-de-La-Libertad.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2017/09/Puerto-de-La-Libertad.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/plaza-marinera-estaria-lista-en-primer-trimestre-de-2019/">Plaza Marinera estaría lista en primer trimestre de 2019</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/cultivar-granos-para-autoconsumo-principal-medio-de-vida-de-los-hogares-vulnerables/">Cultivar granos para autoconsumo, principal medio de vida de los hogares vulnerables</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/hogares-vulnerables-tienden-a-ser-numerosos-y-con-poca-educacion/">Hogares vulnerables tienden a ser numerosos y con poca educación</a></h1>
																															<div class="clear"></div>
					</div>
				</div>
				<!-- -->
				<div class="col-xs-12 col-sm-6 col-md-4">
					<div class="miniBox">
						<h1 class="catName">
							<a href="http://elmundo.sv/category/empresarial">
								EMPRESARIAL
							</a>
						</h1>
						<!-- RECENT POST FROM NACIONALES -->
								
													
														<div class="main-thumbnail">
								<!-- Imagen destacada o primer imagen del post -->
								<a href="http://elmundo.sv/hierromax-de-galvanissa-es-el-acero-de-refuerzo-ideal-para-construccion/" class="thumbnail-wrapper">
								<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Hierromax-construccion-2.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />							
								<!--img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Hierromax-construccion-2.jpg" class="img-responsive thumbnail-wrapper"-->
																</a>

							</div>
							<h1 class="mainPostTitleGlobal"><a href="http://elmundo.sv/hierromax-de-galvanissa-es-el-acero-de-refuerzo-ideal-para-construccion/">Hierromáx de Galvanissa es el acero de refuerzo ideal para construcción</a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/universidad-politecnica-celebro-semana-de-cultura-e-innovacion/">Universidad Politécnica celebró &#8220;Semana de Cultura e Innovación&#8221; </a></h1>
														
															<h1 class="secondPostTitleGlobal"><a href="http://elmundo.sv/jugueton-entrega-donativo-a-plan-internacional/">Juguetón entrega donativo a Plan Internacional</a></h1>
																															<div class="clear"></div>
					</div>
				</div>

				<div class="separador"></div>

			</div>


		</div>
		<div class="col-xs-12 visible-xs visible-sm hidden-md hidden-lg"><hr class="clear"></div>
		<div class="col-xs-12 col-sm-12	col-md-3">	
			
			<div class="col-xs-12 col-sm-6 col-md-12 moreRead nopadding" style="text-align:center;">
				<div class="adblockweb" style="text-align:center;">
	<div id="text-58" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_rect2 -->
<div id='div-gpt-ad-1499235990987-6' style='height:600px; width:300px;'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-6'); });
</script>
</div></div>
		</div></div>			</div>

			<!-- Confidencial -->
			<div class="col-xs-12 col-sm-6 col-md-12 nopadding widget miniBox" style="min-height: 418px!important;">
								<h1 class="MontserratFnt">
					<a href="http://elmundo.sv/category/confidencial">
						CONFIDENCIAL +
					</a>
				</h1>
					
					<div class="customparagraph item1">
						<a href="http://elmundo.sv/confidencial-190318/" class="thumbnail-wrapper">
							<p>Una intensa lucha entre varios sectores del Gobierno y del partido se escenifica desde el …</p>						</a>
					</div>
					
					<div class="customparagraph item2">
						<a href="http://elmundo.sv/confidencial-160318/" class="thumbnail-wrapper">
							<p>Una problemática en la toma de decisiones sobre a quién destituir como funcionario en el …</p>						</a>
					</div>
					
					<div class="customparagraph item3">
						<a href="http://elmundo.sv/confidencial-150318/" class="thumbnail-wrapper">
							<p>Las disputas internas dentro del FMLN están escalando en varias etapas. Dicen que el problema …</p>						</a>
					</div>
							</div>
			<div class="col-xs-12 nopadding widget miniBox" style="min-height:220px!important;">
								<h1 class="MontserratFnt">
					<a href="http://elmundo.sv/category/editorial">
						EDITORIAL +
					</a>
				</h1>
					
					<div class="customPtitle">
						<a href="http://elmundo.sv/la-sociedad-debe-vigilar-la-eleccion-de-la-proxima-sala/" class="thumbnail-wrapper">
							<p>La sociedad debe vigilar la elección de la próxima Sala</p>
						</a>
					</div>
					<div class="parrafoPiquete">
						<p>Los nuevos magistrados deben ser independientes, probos y capaces, sin comp...</p>					</div>
							</div>
			<div class="col-xs-12 hidden-xs visible-sm hidden-md hidden-lg"><hr class="clear"></div>
			<div class="col-xs-12 col-sm-12 col-md-12 nopadding widget miniBox" style="min-height: 395px!important;">
								<h1 class="MontserratFnt">
					<a href="http://elmundo.sv/category/piquete-de-don-mundo">
						PIQUETE DE DON MUNDO +
					</a>
				</h1>
					
										<div class="mainPiquete">
						<a href="http://elmundo.sv/corriendo-hacia-el-abismo/" class="thumbnail-wrapper">
							<p class="lead">Con un bajo crecimiento y excesivo endeudamiento, no hay país que se levante y que salga adelante, el abismo financiero, el fiscal despeñadero y el desastre nacional son su destino final, un gobierno inteligente, responsable y prudente, evita que la &hellip;</p>						</a>
					</div>
										
											<a href="http://elmundo.sv/pagaran-justos-por-pecadores/" class="mostpiquetes">
							Pagarán justos por pecadores						</a>
										
											<a href="http://elmundo.sv/no-nos-quejemos-3/" class="mostpiquetes">
							No nos quejemos						</a>
										
											<a href="http://elmundo.sv/una-gran-responsabilidad/" class="mostpiquetes">
							Una gran responsabilidad						</a>
										
											<a href="http://elmundo.sv/en-que-nos-equivocamos/" class="mostpiquetes">
							¿En qué nos equivocamos?						</a>
												</div>
			
		</div>
	</div>

	<div class="clear separador"></div>

	<div class="row" style="margin-left:0!important; margin-right:0!important;">
		<!-- Post Category Column -->
		<div class="col-xs-12 col-sm-12 col-md-9 nopadding">
			<!-- Google Ads 728x90 -->
		
			<div class="adsense ad728x90">
				 <div class="adblockweb" style="text-align:center;">
	<div id="text-55" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_lead2 -->
<div id='div-gpt-ad-1499235990987-3'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-3'); });
</script>
</div></div>
		</div></div>	
			</div>
		


			
			<!-- Sección para ediciones digitales -->
<h1 class="MontserratFnt" style="color:#000!important;">
	<a href="http://elmundo.sv/category/kiosko-digital/">KIOSKO DIGITAL +</a>
</h1>
<div class="edicionesDigitales">
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
					
				<div class="main-thumbnailDigital">
					<!-- Imagen destacada o primer imagen del post -->
					<a href="http://elmundo.sv/category/e-paper" class="thumbnail-wrapper">
											<img src="http://static.elmundo.sv/kdg-content/featured/mundo/2018/03/mundo190318.jpg" class="img-responsive thumbnail-wrapper" style="width:100%;">
										</a>
				</div>
			</div>
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
					
				<div class="main-thumbnailDigital">
					<!-- Imagen destacada o primer imagen del post -->
					<a href="http://elmundo.sv/category/migueleno" class="thumbnail-wrapper">
											<img src="http://static.elmundo.sv/kdg-content/featured/migueleno/2018/02/migueleno220218.jpg" class="img-responsive thumbnail-wrapper" style="width:100%;">
										</a>
				</div>
			</div>
	<div class="col-xs-12 visible-xs hidden-md hidden-sm"><hr class="clear"></div>
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
		<!-- [+] Periódicos: El Santaneco, Mujer & Familia -->
					
				<div class="main-thumbnailDigital">
					<!-- Imagen destacada o primer imagen del post -->
					<a href="http://elmundo.sv/mujer-familia-28-02-18/" class="thumbnail-wrapper">
											<img src="http://static.elmundo.sv/kdg-content/featured/mujer/2018/02/mujer280218.jpg" class="img-responsive thumbnail-wrapper" style="width:100%;">
										</a>
				</div>
			</div>
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
		<!-- [+] Revistas: VidaSana, Devacaciones, CocinaSana, Bebe & Familia -->
					
				<div class="main-thumbnailDigital">
					<!-- Imagen destacada o primer imagen del post -->
					<a href="http://elmundo.sv/cocina-sana-edicion-4/" class="thumbnail-wrapper">
					<img src="http://static.elmundo.sv/wp-content/uploads/2018/03/Tapa-CocinaSana-04.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />					</a>
				</div>
			</div>
	
			
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
			<div class="main-thumbnailDigital">
				<!-- Imagen destacada o primer imagen del post -->
				<a href="http://elmundo.sv/category/revistas-comerciales" class="thumbnail-wrapper">
				<img src="http://static.elmundo.sv/wp-content/uploads/2017/11/FIAES.jpg" class="img-responsive thumbnail-wrapper wp-post-image" alt="" />				</a>
			</div>
	</div>
	
			
	<div class="col-xs-6 col-sm-2 col-md-2 col-lg-2 noleftpadding">
			<div class="main-thumbnailDigital">
				<!-- Imagen destacada o primer imagen del post -->
				<a href="http://elmundo.sv/category/suplementos-patronales" class="thumbnail-wrapper">
									<img src="http://static.elmundo.sv/kdg-content/featured/suplementos/2018/02/suplementos230218.jpg" class="img-responsive thumbnail-wrapper" style="width:100%;">
								</a>
			</div>
	</div>
		
	<div class="clear"></div>
</div>
<!--div class="col-xs-12">
	<h2 class="secondPostTitleGlobal" style="border-top: 1px solid #eee;padding-top: 10px;">
	<a href="http://elmundo.sv/category/kiosko-digital/">Ver más ediciones digitales</a>
	</h2>
</div-->
			<div class="separador clear"></div>

			
			<!-- Sección para ediciones digitales -->
			<h1 class="MontserratFnt">
				<a href="http://elmundo.sv/category/opinion-grafica">
						OPINIÓN GRÁFICA +
				</a>
			</h1>
			<div>
				<div class="col-xs-12">
											
						<div class="CartoonDEM"><img class="size-full wp-image-881340 aligncenter" src="http://static.elmundo.sv/wp-content/uploads/2018/03/Caricatura-190318.jpg" alt="" />&hellip;</div>
						<p class="fecha" style="font-size: 13px;text-align: center;color: #666;">lunes 19, marzo 2018</p>
									</div>
			</div>

			<div class="separador clear"></div>

		</div>

		<div class="col-xs-12 col-sm-12	col-md-3" id="stickyModul">
			<div class="col-xs-12 nopadding widget">
				<div class="hidden-xs hidden-sm col-md-3 modultop nopadding" style="border-left: 10px solid #ffffff;">
					
					<div class="adblockweb" style="text-align:center;">
	<div id="text-59" class="widget widget_text">			<div class="textwidget"><!-- /12206962/dem_rect3 -->
<div id='div-gpt-ad-1499235990987-7'>
<script>
googletag.cmd.push(function() { googletag.display('div-gpt-ad-1499235990987-7'); });
</script>
</div></div>
		</div></div>					
				</div>
			</div>

			<div class="col-xs-12 nopadding widget miniBox" style="min-height:220px!important;">
								<h1 class="MontserratFnt">
					<a href="http://elmundo.sv/category/buenos-dias">
						BUENOS DÍAS +
					</a>
				</h1>
					
					<div class="customPtitle">
						<a href="http://elmundo.sv/el-nepotismo-cae-mal-y-muy-mal-no-lo-defiendan/" class="thumbnail-wrapper">
							<p>El nepotismo cae mal y muy mal, ¡no lo defiendan!</p>
						</a>
					</div>
					<div class="parrafoPiquete">
						<p>Tristemente hay núcleos familiares enteros enquistados en el Gobierno. Esp...</p>					</div>
							</div>

			<div class="col-xs-12 nopadding widget">
								<h1 class="MontserratFnt">
					<a href="http://elmundo.sv/category/opinion">
						OPINIÓN +
					</a>
				</h1>
					
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/el-plan-de-seguridad-elecciones-2018/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2017/05/Ricardo-Sosa.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Ricardo Sosa</td></tr></table>
							<a href="http://elmundo.sv/el-plan-de-seguridad-elecciones-2018/" class="titleOpinion">
								<p>El plan de seguridad elecciones 2018</p>
							</a>
						</div>
					</div>
																				
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/verguenza-nacional-que-sugiere-cambio/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2016/04/MAURICIO-COLORADO.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Dr. Mauricio Eduardo Colorado</td></tr></table>
							<a href="http://elmundo.sv/verguenza-nacional-que-sugiere-cambio/" class="titleOpinion">
								<p>Vergüenza nacional que sugiere cambio</p>
							</a>
						</div>
					</div>
					<hr class="clear visible-xs visible-sm hidden-md hidden-lg">															
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/peligros-de-la-inminente-alternancia-presidencial/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2016/04/Jorge-Castillo-1.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Jorge Castillo</td></tr></table>
							<a href="http://elmundo.sv/peligros-de-la-inminente-alternancia-presidencial/" class="titleOpinion">
								<p>Peligros de la inminente alternancia presidencial</p>
							</a>
						</div>
					</div>
										<hr class="clear hidden-xs hidden-sm visible-md visible-lg">										
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/factores-que-incidieron-en-el-desplome-del-fmln/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2016/04/jaime-ramirez.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Jaime Ramírez Ortega</td></tr></table>
							<a href="http://elmundo.sv/factores-que-incidieron-en-el-desplome-del-fmln/" class="titleOpinion">
								<p>Factores que incidieron en el desplome del FMLN</p>
							</a>
						</div>
					</div>
															<hr class="clear visible-xs visible-sm hidden-md hidden-lg">					
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/buscando-un-lider/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2016/04/EDUARDO-CALIX.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Eduardo Cálix</td></tr></table>
							<a href="http://elmundo.sv/buscando-un-lider/" class="titleOpinion">
								<p>Buscando un líder</p>
							</a>
						</div>
					</div>
																				
					<div class="col-xs-6 col-sm-6 col-md-4 noleftpadding">
						<div class="main-thumbnail">
							<!-- Imagen destacada o primer imagen del post -->
							<a href="http://elmundo.sv/impulso-oficial-para-el-deporte/" class="thumbnail-wrapper">
							<img src="http://static.elmundo.sv/wp-content/uploads/2016/04/armando-rivera.jpg" class="img-responsive thumbnail-wrapper img-circle wp-post-image" alt="" width="40px" />							</a>

						</div>
						<div>
							<table cellpadding="0" cellspacing="0"><tr><td  class="redactorHome" valign="middle">Armando Rivera Bolaños</td></tr></table>
							<a href="http://elmundo.sv/impulso-oficial-para-el-deporte/" class="titleOpinion">
								<p>Impulso oficial para el deporte</p>
							</a>
						</div>
					</div>
																						</div>
			
		</div>
	</div>
	



<a href="#" title="Ir arriba" class="scrollToTop"><span class="glyphicon glyphicon-chevron-up"></span></a>
<!-- Modal -->
<div class="modal fade bs-example-modal-sm" tabindex="-1" role="dialog" aria-labelledby="mySmallModalLabel">
  <div class="modal-dialog modal-sm" role="document">
    <div class="modal-content">
      <div class="modal-header">
        <button type="button" class="close" data-dismiss="modal" aria-label="Close"><span aria-hidden="true">&times;</span></button>
        <h4 class="modal-title" id="myModalLabel">Formuarlio de búsqueda</h4>
      </div>
      <div class="modal-body">
        <div id="search-2"><form action="http://elmundo.sv/" method="get" class="form-inline" id="busquedadem">

    <fieldset>
		<div class="input-group">
			<input type="text" name="s" id="search" placeholder="Buscar en nuestro sitio web" value="" class="form-control input-sm" />
			<span class="input-group-btn">
				
				<button type="submit" class="btn btn-default btn-sm" id="search_btn"><span class="glyphicon glyphicon-search"></span></button>			
				
			</span>
		</div>
    </fieldset>
</form></div>      </div>
    </div>
  </div>
</div>




<!-- Google Ads 728x90 -->

</div>


<div class="navbar navbar-inverse" style="margin-bottom:0">
	<div class="container">
		<div class="col-xs-12">
			<div class="navbar-header" style="float:none !important;">
				<p class="text-center" style="margin:10px;color:#fff;font-size:12px"><img src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/images/logo-footer.png" width="113" height="23" alt="Diario El Mundo" /><br> Copyright &copy; 2018 Diario El Mundo - Todos los derechos reservados.</p>
			</div>
		</div>
	</div>
</div>



<style>
	.scrollToTop{
		/*width:100px; 
		height:130px;*/
		padding:12px 10px; 
		text-align:center; 
		background: #222;
		font-weight: bold;
		color: #fff;
		text-decoration: none;
		position:fixed;
		bottom:0;
		right:0px;
		display:none;
		z-index: 9999;
		/*background: url('arrow_up.png') no-repeat 0px 20px;*/
	}
	.scrollToTop:hover{
		text-decoration:none;
	}
</style>
<!--[if lt IE 7 ]>
	<script src="//ajax.googleapis.com/ajax/libs/chrome-frame/1.0.3/CFInstall.min.js"></script>
	<script>window.attachEvent('onload',function(){CFInstall.check({mode:'overlay'})});</script>
<![endif]-->	



<script src="https://ajax.googleapis.com/ajax/libs/jquery/1.11.2/jquery.min.js"></script>


<!--div class="popup">
	<h2>EN VIVO | St. Croix Caravelle Hotel & Casino</h2>
	<a class="close" href="#">×</a>
	<div class="content">
		<iframe width="100%" height="200" src="https://www.youtube.com/embed/3Q2CzQclKQc?rel=0&autoplay=1" frameborder="0" allowfullscreen></iframe>
	</div>
</div-->


<script type='text/javascript'>
/* <![CDATA[ */
var countVars = {"disqusShortname":"diarioelmundosv"};
/* ]]> */
</script>
<script type='text/javascript' src='http://elmundo.sv/wp-content/plugins/disqus-comment-system/public/js/comment_count.js?ver=3.0.15'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var pollsL10n = {"ajax_url":"http:\/\/elmundo.sv\/wp-admin\/admin-ajax.php","text_wait":"Tu \u00faltima petici\u00f3n est\u00e1 a\u00fan proces\u00e1ndose. Por favor, espera un momento \u2026","text_valid":"Por favor, elige una respuesta v\u00e1lida para la encuesta.","text_multiple":"N\u00famero m\u00e1ximo de opciones permitidas:","show_loading":"1","show_fading":"1"};
/* ]]> */
</script>
<script type='text/javascript' src='http://elmundo.sv/wp-content/plugins/wp-polls/polls-js.js?ver=2.73.8'></script>
<script type='text/javascript' src='http://cdn.elmundo.sv/wp-includes/js/wp-embed.min.js?ver=4.9.4'></script>





<script>
	jQuery(function(){
		$(".main-menu .menu").addClass("nav navbar-nav");
		$(".main-menu .sub-menu").addClass("dropdown-menu");
		$(".main-menu .menu-item-has-children").each(function(){
			//$(this).removeAttr("class");
			$(this).addClass("dropdown");
			$(this).children().first().addClass("dropdown-toggle");
			//$(this).children().first().attr("data-toggle","dropdown");
		});

	});

	

	$(document).ready(function(){
		//DSQ available content
		$('#comments iframe[title="Disqus"]').hide();


		//--------------------- VIDEO ENVIVO -----------------------
		$(function(){
    		$('.popup').css("visibility", "visible"); 
        	$('.popup').css("opacity", 1); 
        });
  
  		$( ".close" ).click(function() {
	        $('.popup').css("visibility", "hidden"); 
	        $('.popup').css("opacity", 0);
	    });
		//----------------------------------------------------------
		
		//Close Modal
		window.closeModal = function(){
		    $('#emailModal').modal('hide');
		};
		

		//Show menu after webload
					$( "#menu-menu-principal-sin-submenu-2" ).show();
		
		//Check to see if the window is top if not then display button
		$(window).scroll(function(){
			if ($(this).scrollTop() > 100) {
				$(".slicknav_menu").addClass("navbar-fixed-top");
				$('.scrollToTop').fadeIn();
			} else {
				$('.scrollToTop').fadeOut();
				$(".slicknav_menu").removeClass("navbar-fixed-top");
			}
		});
		
		//Click event to scroll to top
		$('.scrollToTop').click(function(){
			$('html, body').animate({scrollTop : 0},800);
			return false;
		});

		//-----------------------------------------------------------
		/* Hamburguer Main menu */
		$( ".cross" ).hide();
		$( ".hamburger" ).hide();
		//$( ".hamburgerMenu" ).hide();
		
		$( ".hamburger" ).click(function() {
			$( "#wrapMenu" ).slideToggle( "fast", function() {
				$( ".hamburger" ).hide();
				$( ".cross" ).show();
				$( "#wrapMenu").show();
				$( ".hamburgerMenu" ).show();
				$( ".sharedNets" ).show();
				$( ".ps__scrollbar-y-rail" ).show();
			});
		});

		$( ".cross" ).click(function() {
			$( "#wrapMenu" ).slideToggle( "fast", function() {
				$( ".cross" ).hide();
				$( ".hamburger" ).show();
				$( "#wrapMenu").hide();
				$( ".hamburgerMenu" ).hide();
				$( ".sharedNets" ).hide();
				$( ".ps__scrollbar-y-rail" ).hide();
			});
		});

		/* Image distribution */
		$(".CartoonDEM img").each(function(){
		    var $this = $(this);
		    if ($this.width() > $this.height()) {
		        $this.addClass("horizontal");
		    }else{
		    	$this.addClass("vertical");
		    }
		});

		//-----------------------------------------------------------
		

			//Sticky navigation nav
			$(window).bind('scroll', function() {
				var navHeight 	= 170; // custom nav height ANTES: 230
				//Put the Mainmenu al the top fixed
				if($(window).scrollTop() > navHeight) {
					$('#menu_principal').addClass('goToTop animated fadeInDown');
					//Ocultamos el menu si esta desplegado y hacemos scrollup
					//$( ".hamburgerMenu" ).hide();
					
					$( ".hamburger" ).show();
					$( ".btnHomepage" ).show();
					$( ".btnSearch" ).show();
					$( ".cross" ).hide();
					$( "#wrapMenu").hide();
					$( ".ps__scrollbar-y-rail" ).hide();

					
					$('#wrapNav').css('display','none');
					$('#imgBrand').css('display', 'block');
					$('#searchBrand').css('display', 'block');
				}else{
					$('#menu_principal').removeClass('goToTop animated fadeInDown');
					//Ocultamos el menu si esta desplegado y hacemos scrollup
					//$( ".hamburgerMenu" ).hide();
					
					$( ".hamburger" ).hide();
					$( ".btnHomepage").hide();
					$( ".btnSearch" ).hide();
					$( ".cross" ).hide();
					$( "#wrapMenu").hide();
					$( ".ps__scrollbar-y-rail" ).hide();
					

					$('#wrapNav').css('display','block');
					$('#imgBrand').css('display', 'none');
					$('#searchBrand').css('display', 'none');
				}

				//LogoMovil DEM
				//($(window).scrollTop() > navHeight) ? setTimeout(function(){ $('#logoFixed').addClass('slideInDown animated noOpacity'); }, 320) : $('#logoFixed').removeClass('slideInDown animated noOpacity');
				//Menu Wordpress
				//($(window).scrollTop() > navHeight) ? $('#NavMainMenu').addClass('fadeInLeft animated') : $('#NavMainMenu').removeClass('fadeInLeft animated');

			});
		


		//Creamos una separacion entre la parte superior del sitio respecto al contenido
		/*$(window).bind('scroll', function() {
			var bheight		= 300; //custom body height
			//Put the Mainmenu al the top fixed
			($(window).scrollTop() > bheight) ? $('body').addClass('MoveContent') : $('body').removeClass('MoveContent');

		});*/
		
		//-----------------------------------------------------------

	});

</script>


<script src="http://cdn.elmundo.sv/wp-content/themes/theme_elmundosv2017/js/perfect-scrollbar.min.js"></script>
<script>
  $(function() {
    Ps.initialize(document.getElementById('wrapMenu'));
  });
</script>
</body>
</html>

<!--
Performance optimized by W3 Total Cache. Learn more: https://www.w3-edge.com/products/

Almacenamiento en caché de objetos 6678/880 objetos que utilizan disk
Page Caching using disk: enhanced 
Red de Entrega de Contenido vía Amazon Web Services: CloudFront: cdn.elmundo.sv
Minificado usando disk
Caching de base de datos 5/104 consultas en 1.066 segundos usando disk

Served from: elmundo.sv @ 2018-03-19 18:22:34 by W3 Total Cache
-->