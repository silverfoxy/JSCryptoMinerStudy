<!DOCTYPE html>
<html lang="es">
<head>
    <meta charset="utf-8">
	<meta http-equiv="content-type" content="text/html; charset=utf-8">
    <meta name="viewport" content="width=device-width, initial-scale=1.0">
    <meta name="description" content="Free business HTML theme fromm ShapeBootstrap, converted for OctoberCMS">
	<meta name="keywords" content="">
    <meta name="author" content="">
    <title>Universidad de El Salvador | Universidad de El Salvador</title>
	
	<!-- core CSS -->
		<link href="http://www2.ues.edu.sv/combine/f5f712950c0c1d1e13a646cc0e8c967b-1508259357" rel="stylesheet">
    <link rel="shortcut icon" href="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ico/favicon.ico">
    <link rel="apple-touch-icon-precomposed" sizes="144x144" href="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ico/144.png">
    <link rel="apple-touch-icon-precomposed" sizes="114x114" href="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ico/114.png">
    <link rel="apple-touch-icon-precomposed" sizes="72x72" href="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ico/72.png">
    <link rel="apple-touch-icon-precomposed" href="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ico/57.png">
</head><!--/head-->

<body class="homepage">

<header id="header">
		<div class="top-bar">
            <div class="container">
                <div class="row">
                        <div class="col-sm-3 col-xs-8">
                            <div class="top-number">
                                <p><i class="fa fa-phone-square"></i> +(503)2511-2000</p>
                            </div>
                        </div>
                        

                        
                        <div class="col-sm-3 col-xs-8">
                                <div class="social">
                                      <ul class="social-share">
                                          <li><a href="https://www.facebook.com/UESoficial.SV/"><i class="fa fa-facebook"></i></a></li>
                                          <li><a href="https://twitter.com/UESoficial"><i class="fa fa-twitter"></i></a></li>
                                          <li><a href="http://www.ues.edu.sv/rss.xml"><i class="fa fa-rss"></i></a></li> 
                                          <li><a href="http://www.ues.edu.sv/rss.xml"><i class="fa fa-whatsapp"></i></a></li> 
                                       </ul>
                                </div>
                        </div>
                                                <div class="col-sm-6 col-xs-8">
                                <nav class="navbar2 top-nav">
  <div class="container-fluid">
    <div class="navbar-header">
      <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#myNavbar">
        <span class="icon-bar"></span>
        <span class="icon-bar"></span>
        <span class="icon-bar"></span>
      </button>

    </div>
    <div class="collapse navbar-collapse" id="myNavbar">
      <ul class="navbar2 top-nav">
        <li><a href="nuestra-universidad">Nuestra Universidad     </a></li>
        <li><a href="administracion">Administración     </a></li>
        <li><a href="http://www.transparencia.ues.edu.sv/">Portal de Transparencia</a></li>
      </ul>
    </div>
  </div>
</nav>                        </div>
                </div><!--/.row-->
            </div><!--/.container-->
	</div><!--/.top-bar-->        



<nav class="navbar navbar-inverse" role="banner">
	<div class="container">
		<div class="navbar-header">
			<button type="button" class="navbar-toggle" data-toggle="collapse" data-target=".navbar-collapse">
			<span class="sr-only">Toggle navigation</span>
			<span class="icon-bar"></span>
			<span class="icon-bar"></span>
			<span class="icon-bar"></span>
			</button>
			<a class="navbar-brand" href=""><img src="http://www2.ues.edu.sv/themes/UES-THEME/assets/images/ues_logo3.svg" alt="logo"></a>
	<div id="header_front"><h1 style="color:#fff">Universidad de El Salvador</h1><h4 style="color:#fff">"HACIA LA LIBERTAD POR LA CULTURA"</h4></div></div>
		<div class="collapse navbar-collapse">
			<ul class="nav navbar-nav navbar-right">
				            <li class=" ">
            <a href="http://www2.ues.edu.sv"
                                class="">
                Inicio
                            </a>
                    </li>
            <li class=" ">
            <a href="http://www2.ues.edu.sv/estudiantes"
                                class="">
                Estudiantes
                            </a>
                    </li>
            <li class=" ">
            <a href="http://www2.ues.edu.sv/facultades"
                                class="">
                Facultades
                            </a>
                    </li>
            <li class=" ">
            <a href="http://www2.ues.edu.sv/proyeccion-social"
                                class="">
                Proyección Social
                            </a>
                    </li>
            <li class=" ">
            <a href="http://www2.ues.edu.sv/investigacion"
                                class="">
                Investigación
                            </a>
                    </li>
    
			</ul>
			
		</div>
	</div>
</nav><!--/nav-->  

</header><!--/header-->

    <section id="carousel portal">
    <div class="container">	
    
     <div id="front_slide" class="carousel slide" data-ride="carousel">
  <!-- Indicators -->
  <ol class="carousel-indicators">
    <li data-target="front_slide" data-slide-to="0" class="active"></li>
    <li data-target="front_slide"data-slide-to="1"></li>
    <li data-target="front_slide" data-slide-to="2"></li>
    <li data-target="front_slide" data-slide-to="3"></li>
  </ol>

  <!-- Wrapper for slides -->
  <div class="carousel-inner" role="listbox">
    <div class="item active"> 
      <img class="img-responsive" src="http://www.ues.edu.sv/storage/app/media/Carousel_img3/Residuos de Cafe.jpg" alt="analisis">

    </div>

    <div class="item">
      <img class="img-responsive" src="http://www.ues.edu.sv/storage/app/media/Carousel_img3/Salud Sexual-.jpg" alt="salud sexual">
    </div>



  </div>

  <!-- Left and right controls -->
  <a class="left carousel-control" href="#front_slide" role="button" data-slide="prev">
    <span class="glyphicon glyphicon-chevron-left" aria-hidden="true"></span>
    <span class="sr-only">Previous</span>
  </a>
  <a class="right carousel-control" href="#front_slide" role="button" data-slide="next">
    <span class="glyphicon glyphicon-chevron-right" aria-hidden="true"></span>
    <span class="sr-only">Next</span>
  </a>
</div>     <!--   <a class="prev hidden-xs" href="#main-slider" data-slide="prev">
        <i class="fa fa-chevron-left"></i>
        </a>
        <a class="next hidden-xs" href="#main-slider" data-slide="next">
        <i class="fa fa-chevron-right"></i>
        </a>-->
     </div>
</section>




<section id="noticias">
    <div class="container">	
          <div class="col-sm-4 wow fadeInDown">

             
      <div class="feature-wrap"><i class="fa fa-bullhorn"></i><h3>Cartelera</h3></div>
      <div class="well"><a href="http://www.ues.edu.sv/storage/app/media/avisos/pronunciamientoUES.jpg"><img class="img-responsive"  src="http://www.ues.edu.sv/storage/app/media/avisos/pronunciamientoUES.jpg" alt="pronunciamiento"></a>
             </div>
             
     <div class="well"><a href="http://distancia.ues.edu.sv/"><img class="img-responsive"  src="http://www.ues.edu.sv/storage/app/media/avisos/adistancia.png" alt="Educacion a distancia"> </a></div>

                   <!-- <div class="well"><a href="http://www.ues.edu.sv/storage/app/media/avisos/acuedo-n-003-2017-2019-viii-62.jpg"><img class="img-responsive"  src="http://www.ues.edu.sv/storage/app/media/avisos/acuedo-n-003-2017-2019-viii-62.jpg" alt="foro juventud"> </a>
             </div>
                  
                  
                  
                  <div class="well"><a href="  http://www.ues.edu.sv/storage/app/media/Documentos/Rendicion_de_Cuentas_2016.pdf">Rendición de Cuentas</a>
             </div>
                 <div class="well"><a href="http://www.ues.edu.sv/storage/app/media/avisos/ciencias_forenses.jpg"><img class="img-responsive"  src="http://www.ues.edu.sv/storage/app/media/avisos/ciencias_forenses.jpg" alt="ciencias_forenses"> </a>
             </div>
            
                 <div class="well"><a href="  http://www.ues.edu.sv/storage/app/media/Documentos/Los_Cobanos_tortugas_informe.pdf">Informe Técnico.
Evento de mortandad de tortugas marinas</a>
             </div>

          

              <div class="well"><a href="http://www.ues.edu.sv/storage/app/media/uploaded-files/doc03575520170815145822.pdf"><h4>Dirección General de Protección Civil, Prevención y Mitigación de Desastres</h4></br>
Resultados de la evaluación de infraestructura de los edificios que resultaron dañados en el marco de la alerta amarilla decretada por el sismo de 5.1 del 10 de abril de 2017.
</a>
             </div>    <div class="well"><a href="http://www.ues.edu.sv/storage/app/media/uploaded-files/doc03575720170815150156.pdf"><h4>Desarrollo Físico de la UES presentó informe al CSU </h4></br>
Reporte preliminar de evaluación de daños de infraestructura del campus, causado por el enjambre sísmico en el periodo comprendido entre el 9 y 10 de abril. 

</a>
             </div>-->
             
             
  
             <!--<div class="well"><h4>Aviso</h4> 
A los graduandos se les comunica que para cualquier información sobre las graduaciones consultar el sitio de la Secretaría de Asuntos Académicos: <a href="http://saa.ues.edu.sv/portal">http://saa.ues.edu.sv/portal</a>
             </div> -->
              
                        
 
</div>   <div class="col-sm-4">
                                
        <div class="cartelera">
            <div class="well">  
                  <div class="text-center"> <h3>8 de marzo</h3><h4> Día Internacional de la Mujer</h4>
                    <p><a href="storage/app/media/avisos/mujer dia.jpg"><img class="img-responsive" src="storage/app/media/avisos/mujer dia.jpg" alt="mujer"></a></p>
                </div>
            </div>
            <div class="well">   
                    <iframe width="" height="" src="https://www.youtube.com/embed/CzF6SwrTFCs" frameborder="0" allow="autoplay; encrypted-media" allowfullscreen></iframe>
            </div>

        </div>
        
</div>  
       <div class="col-sm-4 wow fadeInDown">

    <div class="indice">    
        <div class="panel panel-default">
            <div class="panel-body">
                <div class="feature-wrap">
                    <i class="fa fa-search"></i><h4>Búsqueda</h4>
                </div>

                <div class="search">
                           <form action="http://www2.ues.edu.sv/search" method="get">
    <input name="q" type="text" placeholder="búsqueda" autocomplete="off">
    <button type="submit">Buscar</button>
</form> 
                </div>
                </div>
                

            <div class="panel-body">
                <div class="feature-wrap">
                    <i class="fa fa-phone"></i><h4>Directorio </h4>
                         <p>Conmutador UES: 2511-2000</p>
                      <a href="directorio"><p>Enlace a Oficinas Centrales</p></a>
                </div>
            </div>
        
        <div class="panel-body">
            <div class="feature-wrap">
                    <a href="https://correo.ues.edu.sv/login/module.php/core/loginuserpass.php?AuthState=_11ba3a856a215cc0683961963fda1400e3f91dfce5%3Ahttps%3A%2F%2Fcorreo.ues.edu.sv%2Flogin%2Fsaml2%2Fidp%2FSSOService.php%3Fspentityid%3Dgoogle.com%26cookieTime%3D1487692519%26RelayState%3Dhttps%253A%252F%252Fwww.google.com%252Fa%252Fues.edu.sv%252FServiceLogin%253Fservice%253Dmail%2526passive%253Dtrue%2526rm%253Dfalse%2526continue%253Dhttps%25253A%25252F%25252Fmail.google.com%25252Fmail%25252F%2526ss%253D1%2526ltmpl%253Ddefault%2526ltmplcache%253D2%2526emr%253D1%2526osid%253D1"><i class="fa fa-envelope-o"></i><h4>Correo Electrónico Institucional UES </h4></a>
                    <!--<p>Correo Electrónico Institucional de la Universidad de El Salvador</p>-->
            </div>
        </div>
        
                <div class="panel-body">
            <div class="feature-wrap">
                    <a href="medios"><i class="fa fa-camera"></i><h4>Medios Universitarios</h4></a>
                    <p></p>
            </div>
        </div>
        
    </div>  </div>

</div>       
     </div>
</section>
<!--<section id="medios">    
      <div class="center wow fadeInDown">
          <h1>Medios Universitarios</h1>
       </div>
     <div class="container">
       <div class="row">
     Aqui se puede colocar el partial "medios"
       
       
       </div>
     </div>
</section> -->
<!--<section id="medios">
    <div class="container">	
  
     </div>
</section>-->
<section id="bottom">
<div class="container wow fadeInDown" data-wow-duration="1000ms" data-wow-delay="600ms">
        <div class="row">
            <div class="col-md-3 col-sm-6">
                <div class="widget">
                 <h3>Secretarias</h3>
                    <ul class="list-group">  
                        <li><a href="http://secretariageneral.ues.edu.sv/">Secretaría General</a></li>
                       <li><a href="http://saa.ues.edu.sv/portal/">Secretaría de Asuntos Académicos</a></li>
                         <li><a href="http://proyeccionsocial.ues.edu.sv/">Secretaría de Proyección Social</a></li>
                     <li><a href="http://www.eluniversitario.ues.edu.sv/">Secretaría de Comunicaciones</a></li>
                      <li><a href="https://es-es.facebook.com/ArteyCulturaUES/">Secretaría de Arte y Cultura</a></li>
                         <li><a href="http://www.bienestar.ues.edu.sv/">Secretaría de Bienestar Universitario</a></li>
                        <li><a href="http://www.ues.edu.sv/secretaria-de-relaciones-nacionales-e-internacionales/">Secretaría de Relaciones</a></li>
                         <li><a href="en-construccion">Secretaría de Planificación</a></li>
                    </ul> 
                </div>    
            </div><!--/.col-md-3-->

           
            <div class="col-md-3 col-sm-6">
                <div class="widget">
                    <h3>Contactos</h3>
                     <ul>
                        <li><a href="http://www.csuca.org/">Consejo Superior Centroamericano</a></li>
                   
    
                        <li><a href="programa-de-graduados">Programa de Estudios de Graduados</a></li>
                    <!--         <li><a href=">Consejo Centroamericano de Acreditación de la Educación Superior</a></li>-->
                        <li><a href="http://redgira.unanleon.edu.ni/organizacion.html">Red Gira</a></li>
                        <li><a href="http://cca.ucr.ac.cr/">Consejo Centroamericano de Acreditación de la Educación Superior</a></li>
                    </ul> 
                </div>    
            </div><!--/.col-md-3-->

            <div class="col-md-3 col-sm-6">
                <div class="widget">
                    <h3>Indicadores</h3>
                    <ul>
                        <li><a href="#">Inicio</a></li>
                        <li><a href="indicadores">Derechos Reservados</a></li>
                        <li><a href="en-construccion">Mapa del Sitio</a></li>
                        <li><a href="indicadores">Contacto UES </a></li> 
                    </ul>
                </div>    
            </div><!--/.col-md-3-->

            <div class="col-md-3 col-sm-6">
                <div class="widget">
                    <h3>Servicios</h3>
                    <ul>
						<li><a href="http://biblioteca.ues.edu.sv/portal/">Sistema Bibliotecario</a></li>
						<li><a href="http://www.ues.edu.sv/unidad_calidad/">Unidad Técnica de Gestión de la Calidad</a></li>
						<li><a href="http://www.editorialuniversitaria.ues.edu.sv/">Editorial Universitaria</a></li>
                        <li><a href="http://www.ues.edu.sv/libreria/">Librería Universitaria</a></li>
                        <li><a href="https://www.facebook.com/pages/CENIUES/">CENIUES</a></li>
                        <li><a href="http://www.ues.edu.sv/fup/">Fondo Universitario de Protección</a></li>
                    </ul>
                </div>    
            </div><!--/.col-md-3-->
        </div>
    </div><section><!--/#bottom-->

<footer id="footer" class="midnight-blue">
	<div class="container">
        <div class="row">
            <div class="col-sm-7">
				&copy;  2018 Universidad de El Salvador. Todos los derechos reservados.</br> Ciudad Universitaria, Final de Av.Mártires y Héroes del 30 julio, San Salvador, El Salvador, América Central. Teléfonos: +(503) 2511-2000 
            </div>
            <div class="col-sm-5">
                <ul class="pull-right">
                       <li><a href="#">Inicio</a></li>
                        <li><a href="indicadores">Derechos Reservados</a></li>
                        <li><a href="en-construccion">Mapa del Sitio</a></li>
                        <li><a href="indicadores">Contacto UES </a></li> 
                </ul>
            </div>
        </div>
    </div>
    

<!-- Piwik -->
<script type="text/javascript">
  var _paq = _paq || [];
  // tracker methods like "setCustomDimension" should be called before "trackPageView"
  _paq.push(['trackPageView']);
  _paq.push(['enableLinkTracking']);
  (function() {
    var u="//www.ues.edu.sv/webanalisis/";
    _paq.push(['setTrackerUrl', u+'piwik.php']);
    _paq.push(['setSiteId', '1']);
    var d=document, g=d.createElement('script'), s=d.getElementsByTagName('script')[0];
    g.type='text/javascript'; g.async=true; g.defer=true; g.src=u+'piwik.js'; s.parentNode.insertBefore(g,s);
  })();
</script>
<!-- End Piwik Code --></footer><!--/#footer-->

<!-- Scripts -->
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/html5shiv.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/respond.min.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/jquery.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/bootstrap.min.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/jquery.prettyPhoto.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/jquery.isotope.min.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/main.js"></script>
<script type="text/javascript" src="http://www2.ues.edu.sv/themes/UES-THEME/assets/js/wow.min.js"></script>
<script src="/modules/system/assets/js/framework.js"></script>
<script src="/modules/system/assets/js/framework.extras.js"></script>
<link rel="stylesheet" property="stylesheet" href="/modules/system/assets/css/framework.extras.css">
             
                           

<!-- Piwik -->
<script type="text/javascript">
  var _paq = _paq || [];
  // tracker methods like "setCustomDimension" should be called before "trackPageView"
  _paq.push(['trackPageView']);
  _paq.push(['enableLinkTracking']);
  (function() {
    var u="//www.ues.edu.sv/webanalisis/";
    _paq.push(['setTrackerUrl', u+'piwik.php']);
    _paq.push(['setSiteId', '1']);
    var d=document, g=d.createElement('script'), s=d.getElementsByTagName('script')[0];
    g.type='text/javascript'; g.async=true; g.defer=true; g.src=u+'piwik.js'; s.parentNode.insertBefore(g,s);
  })();
</script>
<!-- End Piwik Code -->


</body>
</html>