<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML 1.0 Transitional//EN" "http://www.w3.org/TR/xhtml1/DTD/xhtml1-transitional.dtd"> <html xmlns="http://www.w3.org/1999/xhtml">
<head>

<script language="JavaScript" src="js/jquery-1.10.2.js"></script>
<script language="JavaScript" src="js/jquery-ui/jquery-ui.js"></script>
<script language="JavaScript" src="js/jquery-browser.js"></script>
<script language="JavaScript" src="js/jquery.form.js"></script>

<script language="JavaScript" src="js/js2013.js"></script>

<link href="css/style2.css" type="text/css" rel="stylesheet">
<link href="js/jquery-ui/jquery-ui.min.css" type="text/css" rel="stylesheet">

<link rel="shortcut icon" href="img/favicon.png" />

<meta http-equiv="Content-Type" content="text/html; charset=utf-8" />
<meta name="Keywords" content="Universidad,Francisco,Gavidia,">
<meta name="Description" content="Universidad Francisco Gavidia">

<title>::Universidad Francisco Gavidia::</title>
<script language="JavaScript">
(function(a){jQuery.browser.mobile=/android.+mobile|avantgo|bada/|blackberry|blazer|compal|elaine|fennec|hiptop|iemobile|ip(hone|od)|iris|kindle|lge |maemo|midp|mmp|netfront|opera m(ob|in)i|palm( os)?|phone|p(ixi|re)/|plucker|pocket|psp|symbian|treo|up.(browser|link)|vodafone|wap|windows (ce|phone)|xda|xiino/i.test(a)||/1207|6310|6590|3gso|4thp|50[1-6]i|770s|802s|a wa|abac|ac(er|oo|s-)|ai(ko|rn)|al(av|ca|co)|amoi|an(ex|ny|yw)|aptu|ar(ch|go)|as(te|us)|attw|au(di|-m|r |s )|avan|be(ck|ll|nq)|bi(lb|rd)|bl(ac|az)|br(e|v)w|bumb|bw-(n|u)|c55/|capi|ccwa|cdm-|cell|chtm|cldc|cmd-|co(mp|nd)|craw|da(it|ll|ng)|dbte|dc-s|devi|dica|dmob|do(c|p)o|ds(12|-d)|el(49|ai)|em(l2|ul)|er(ic|k0)|esl8|ez([4-7]0|os|wa|ze)|fetc|fly(-|_)|g1 u|g560|gene|gf-5|g-mo|go(.w|od)|gr(ad|un)|haie|hcit|hd-(m|p|t)|hei-|hi(pt|ta)|hp( i|ip)|hs-c|ht(c(-| |_|a|g|p|s|t)|tp)|hu(aw|tc)|i-(20|go|ma)|i230|iac( |-|/)|ibro|idea|ig01|ikom|im1k|inno|ipaq|iris|ja(t|v)a|jbro|jemu|jigs|kddi|keji|kgt( |/)|klon|kpt |kwc-|kyo(c|k)|le(no|xi)|lg( g|/(k|l|u)|50|54|e-|e/|-[a-w])|libw|lynx|m1-w|m3ga|m50/|ma(te|ui|xo)|mc(01|21|ca)|m-cr|me(di|rc|ri)|mi(o8|oa|ts)|mmef|mo(01|02|bi|de|do|t(-| |o|v)|zz)|mt(50|p1|v )|mwbp|mywa|n10[0-2]|n20[2-3]|n30(0|2)|n50(0|2|5)|n7(0(0|1)|10)|ne((c|m)-|on|tf|wf|wg|wt)|nok(6|i)|nzph|o2im|op(ti|wv)|oran|owg1|p800|pan(a|d|t)|pdxg|pg(13|-([1-8]|c))|phil|pire|pl(ay|uc)|pn-2|po(ck|rt|se)|prox|psio|pt-g|qa-a|qc(07|12|21|32|60|-[2-7]|i-)|qtek|r380|r600|raks|rim9|ro(ve|zo)|s55/|sa(ge|ma|mm|ms|ny|va)|sc(01|h-|oo|p-)|sdk/|se(c(-|0|1)|47|mc|nd|ri)|sgh-|shar|sie(-|m)|sk-0|sl(45|id)|sm(al|ar|b3|it|t5)|so(ft|ny)|sp(01|h-|v-|v )|sy(01|mb)|t2(18|50)|t6(00|10|18)|ta(gt|lk)|tcl-|tdg-|tel(i|m)|tim-|t-mo|to(pl|sh)|ts(70|m-|m3|m5)|tx-9|up(.b|g1|si)|utst|v400|v750|veri|vi(rg|te)|vk(40|5[0-3]|-v)|vm40|voda|vulc|vx(52|53|60|61|70|80|81|83|85|98)|w3c(-| )|webc|whit|wi(g |nc|nw)|wmlb|wonu|x700|xda(-|2|g)|yas-|your|zeto|zte-/i.test(a.substr(0,4))})(navigator.userAgent||navigator.vendor||window.opera);

function setCookie(cname,cvalue,exdays)
{
var d = new Date();
d.setTime(d.getTime()+(exdays*24*60*60*1000));
var expires = "expires="+d.toGMTString();
document.cookie = cname + "=" + cvalue + "; " + expires;
}

function getCookie(cname)
{
var name = cname + "=";
var ca = document.cookie.split(';');
for(var i=0; i<ca.length; i++)
{
var c = ca[i].trim();
if (c.indexOf(name)==0) return c.substring(name.length,c.length);
}
return "";
}

var medio='';
var cMedio=getCookie('medio');
if (cMedio.length>0) {medio=cMedio;}

var parametros = {};
location.search.substr(1).split("&").forEach(function(item) {parametros[item.split("=")[0]] = item.split("=")[1]})
if (parametros['medio']) {medio=parametros['medio'];}
setCookie('medio',medio,365);

if ((jQuery.browser.mobile && medio=='') || medio=='movil') {
window.location = "http://www.ufg.edu.sv/m.index.html";
}
</script>
<style type="text/css">
<!--
body {
margin-left: 0px;
margin-top: 0px;
margin-right: 0px;
margin-bottom: 0px;
background-image: url(img/fondo2.jpg);
background-repeat: repeat-x;
}
-->
</style>

<style type="text/css">
<!--
#apDiv1 {
position:absolute;
left:41px;
top:4px;
width:1019px;
height:671px;
z-index:1;
}
#apDiv2 {
position: absolute;
margin-left: 210px;
top:0px;
width:927px;
height:800px;
z-index:1;
background-color: #99FF00;
}
#apDiv3 {
position:absolute;
left: 50%;
margin-left: -464px;
top:0px;
width:927px;
height:1500px;
z-index:1;
}
#apDiv4 {
position:absolute;
left:0px;
top:0px;
width:927px;
height:136px;
z-index:0;
}
#apDiv5 {
position:absolute;
left:0px;
top:137px;
width:205px;
height:760px;
z-index:3;
}
#apDiv6 {
position:absolute;
left:217px;
top:137px;
width:710px;
height:798px;
z-index:2;
}
#apDiv7 {
position:absolute;
left:0px;
/*top:1005px;*/
top:1020px;
width:927px;
height:95px;
z-index:2;
font-size:
}
#apDiv8 {
position:absolute;
left:0px;
top:4px;
width:637px;
height:75px;
z-index:2;
}
#apDiv9 {
position:absolute;
left:722px;
top:42px;
width:185px;
height:29px;
z-index:2;
}
#apDiv10 {
position:absolute;
left:728px;
top:21px;
width:162px;
height:20px;
z-index:2;
background-color: #FFFFFF;
}
#apDiv11 {
position:absolute;
left:895px;
top:21px;
width:25px;
height:20px;
z-index:2;
}
#apDiv12 {
position:absolute;
left:720px;
top:2px;
width:209px;
height:18px;
z-index:2;
}
#apDiv13 {
position:absolute;
left:0px;
top:83px;
width:927px;
height:3px;
z-index:2;
background-color: #FF6600;
}
#apDiv14 {
position:absolute;
left:0px;
top:97px;
width:927px;
height:28px;
z-index:2;
}
#apDiv15 {
position:absolute;
left:0px;
top:0px;
width:710px;
height:329px;
z-index:2;

}
#apDiv16 {
position:absolute;
left:0px;
top:330px;
width:710px;
height:15px;
z-index:2;
vertical-align: middle;
}
#apDiv17 {
position:absolute;
left:0px;
top:10px;
width:569px;
height:20px;
z-index:2;
}
#apDiv18 {
position:absolute;
left:0px;
top:475px;
width:927px;
height:3px;
z-index:2;
background-color: #0066FF;
}
#apDiv19 {
position:absolute;
left:0px;
top:0px;
width:205px;
height:327px;
z-index:2;
background-image: url(img/fondo-menu-izq.jpg);
border-color: #00CCFF;
border-width: 1px;
border-style: solid;
border-radius:0px;
-moz-border-radius:0px; /* Firefox */
-webkit-border-radius:0px; /* Safari y Chrome */
}
#apDiv20 {
position:absolute;
left:0px;
top:351px;
width:205px;
height:54px;
z-index:2;
}
#apDiv21 {
position:absolute;
left:0px;
top:469px;
width:205px;
height:54px;
z-index:2;
}
#apDiv22 {
position:absolute;
left:0px;
/*top:587px;*/
top:647px;
width:203px;
/*height:239px;*/
height:209px;
z-index:2;
overflow: auto;
border-color: #004B97;
border-width: 1px;
border-style: solid;
border-radius:0px;
-moz-border-radius:0px; /* Firefox */
-webkit-border-radius:0px; /* Safari y Chrome */
}
#apDiv23 {
position:absolute;
left:0px;
top:665px;
width:708px;
height:95px;
z-index:2;
border-color: #004B97;
border-width: 1px;
border-style: solid;
border-radius:6px;
-moz-border-radius:6px; /* Firefox */
-webkit-border-radius:6px; /* Safari y Chrome */
}
#apDiv24 {
position:absolute;
left:0px;
top:4px;
width:708px;
height:86px;
z-index:2;
}
#apDiv25 {
position:absolute;
left:5px;
top:9px;
width:193px;
height:62px;
z-index:2;
}
#apDiv26 {
position:absolute;
left:5px;
top:79px;
width:193px;
height:88px;
z-index:2;
}
#apDiv27 {
position:absolute;
left:80px;
top:175px;
width:46px;
height:16px;
z-index:2;
}

#apDiv28 {
position:absolute;
left:0px;
top:375px;
width:440px;
height:453px;
z-index:2;
}
#apDiv29 {
position:absolute;
left:450px;
top:375px;
width:260px;
/*height:453px;*/
height:485px;
z-index:2;
}
#apDiv30 {
position:absolute;
left:445px;
top:376px;
width:1px;
/*height:450px;*/
height:490px;
z-index:2;
background-color: #004B97;
}

#apDiv31 {
position:absolute;
left:516px;
top:302px;
width:158px;
height:14px;
z-index:2;
}
#apDiv32 {
position:absolute;
left:0px;
top:3px;
width:13px;
height:12px;
z-index:2;
}
#apDiv33 {
position:absolute;
left:22px;
top:1px;
width:14px;
height:14px;
z-index:2;
border-top: 1px solid #ffffff;
border-right: 1px solid #ffffff;
border-bottom: 1px solid #ffffff;
border-left: 1px solid #ffffff;
}
#apDiv34 {
position:absolute;
left:45px;
top:1px;
width:14px;
height:14px;
z-index:3;
border-top: 1px solid #ffffff;
border-right: 1px solid #ffffff;
border-bottom: 1px solid #ffffff;
border-left: 1px solid #ffffff;
}
#apDiv35 {
position:absolute;
left:69px;
top:1px;
width:14px;
height:14px;
z-index:4;
border-top: 1px solid #ffffff;
border-right: 1px solid #ffffff;
border-bottom: 1px solid #ffffff;
border-left: 1px solid #ffffff;
}
#apDiv36 {
position:absolute;
left:94px;
top:1px;
width:14px;
height:14px;
z-index:5;
border-top: 1px solid #ffffff;
border-right: 1px solid #ffffff;
border-bottom: 1px solid #ffffff;
border-left: 1px solid #ffffff;
}
#apDiv37 {
position:absolute;
left:118px;
top:1px;
width:14px;
height:14px;
z-index:6;
border-top: 1px solid #ffffff;
border-right: 1px solid #ffffff;
border-bottom: 1px solid #ffffff;
border-left: 1px solid #ffffff;
}
#apDiv38 {
position:absolute;
left:166px;
top:3px;
width:13px;
height:11px;
z-index:7;
}
#apDiv39 {
position:absolute;
left:28px;
top:4px;
width:200px;
height:22px;
z-index:2;
}
#apDiv40 {
position:absolute;
left:0px;
top:39px;
width:260px;
/*height:410px;*/
height:445px;
z-index:2;
overflow: scroll;
overflow-x: hidden;
}
#apDiv41 {
position:absolute;
left:145px;
/*top:455px;*/
top:490px;
width:100px;
height:18px;
z-index:2;
}
#apDiv42 {
position:absolute;
left:120px;
top:4px;
width:380px;
height:22px;
z-index:2;
}
#apDiv43 {
position:absolute;
left:20px;
top:39px;
width:400px;
height:245px;
z-index:2;
}
#apDiv44 {
position:absolute;
left:12px;
top:319px;
width:415px;
height:55;
z-index:2;
border-color: #004B97;
border-width: 1px;
border-style: dashed;
overflow: hidden;
}

#apDiv45 {
position:absolute;
left:99px;
top:295px;
width:230px;
height:16px;
z-index:2;
}
#apDiv46 {
position:absolute;
left:0px;
top:3px;
width:13px;
height:12px;
z-index:2;
}
#apDiv47 {
position:absolute;
left:22px;
top:0px;
width:14px;
height:14px;
z-index:3;
}
#apDiv48 {
position:absolute;
left:50px;
top:0px;
width:14px;
height:14px;
z-index:4;
}
#apDiv49 {
position:absolute;
left:78px;
top:0px;
width:14px;
height:14px;
z-index:5;
}
#apDiv50 {
position:absolute;
left:106px;
top:0px;
width:14px;
height:14px;
z-index:6;
}
#apDiv51 {
position:absolute;
left:134px;
top:0px;
width:14px;
height:14px;
z-index:7;
background-color: #FF3300;
}
#apDiv52 {
position:absolute;
left:162px;
top:0px;
width:14px;
height:14px;
z-index:8;
}
#apDiv53 {
position:absolute;
left:190px;
top:0px;
width:14px;
height:14px;
z-index:9;
}
#apDiv54 {
position:absolute;
left:216px;
top:2px;
width:13px;
height:12px;
z-index:10;
}
#apDiv55 {
position:absolute;
left:12px;
top:375px;
/*top:490px;*/
width:415px;
height:55px;
z-index:2;
}
#apDiv56 {
position:absolute;
left:326px;
/*top:455px;*/
top:490px;
width:100px;
height:18px;
z-index:2;
}

#apDiv57 {
position:absolute;
left:0px;
top:410px;
width:205px;
height:54px;
z-index:2;
}
#apDiv58 {
position:absolute;
left:259px;
top:0px;
width:451px;
height:325px;
z-index:2;
border-color: #00CCFF;
border-width: 1px;
border-style: solid;
border-radius:12px;
-moz-border-radius:12px; /* Firefox */
-webkit-border-radius:12px; /* Safari y Chrome */
}
#apDiv59 {
position:absolute;
left:0px;
top:0px;
width:254px;
height:160px;
z-index:2;
border-color: #00CCFF;
border-width: 1px;
border-style: solid;
border-radius:12px;
-moz-border-radius:12px; /* Firefox */
-webkit-border-radius:12px; /* Safari y Chrome */
}
#apDiv60 {
position:absolute;
left:0px;
top:165px;
width:254px;
height:160px;
z-index:2;
border-color: #00CCFF;
border-width: 1px;
border-style: solid;
border-radius:12px;
-moz-border-radius:12px; /* Firefox */
-webkit-border-radius:12px; /* Safari y Chrome */
}
#apDiv61 {
position:absolute;
left:0px;
top:1186px;
width:927px;
height:8px;
z-index:2;
background-color: #004B97;
}

#apDiv78 {
position:absolute;
left:0px;
top:1200px;
width:925px;
height:245px;
z-index:2;
border-color: #004B97;
border-width: 1px;
border-style: solid;
border-radius:1px;
-moz-border-radius:1px; /* Firefox */
-webkit-border-radius:1px;
}
#apDiv79 {
position:absolute;
left:0px;
top:26px;
width:925px;
height:1px;
z-index:2;
background-color: #004b97;
}
#apDiv80 {
position:absolute;
left:13px;
top:-22px;
width:40px;
height:19px;
z-index:2;
}

#apDiv82 {
position:absolute;
left:177px;
top:38px;
width:150px;
height:180;
z-index:2;
line-height: 10px;
}

#apDiv83 {
position:absolute;
left:357px;
top:38px;
width:165px;
height:180;
z-index:2;
}
#apDiv84 {
position:absolute;
left:740px;
top:38px;
width:170px;
height:198px;
z-index:2;
}
#apDiv85 {
position:absolute;
left:547px;
top:38px;
width:165px;
height:183;
z-index:2;
}
#apDiv86 {
position:absolute;
left:18px;
top:38px;
width:130px;
height:180;
z-index:2;
}

#apDiv74 {
position:absolute;
left:0px;
top:587px;
width:205px;
height:55px;
z-index:2;
}

a:link {
text-decoration: none;
}
a:visited {
text-decoration: none;
}
a:hover {
text-decoration: none;
color: #FF3300;
}
a:active {
text-decoration: none;
}

#apDiv62 {
position:absolute;
left:0px;
top:528px;
width:205px;
height:55px;
z-index:2;
}
.style1 {
color: #FFFFFF;
font-weight: bold;
}
#apDiv63 {
position:absolute;
left:822px;
top:1379px;
width:185px;
height:9px;
z-index:2;
}
#apDiv64 {
position:absolute;
left:636px;
top:1378px;
width:185px;
height:9px;
z-index:3;
}
#apDiv65 {
position:absolute;
left:23px;
top:301px;
width:193px;
height:18px;
z-index:2;
}
#apDiv66 {
position:absolute;
left:317px;
top:437px;
width:18px;
height:20px;
z-index:2;
}
#apDiv67 {
position:absolute;
left:27px;
top:0px;
width:16px;
height:16px;
z-index:3;
}
#apDiv68 {
position:absolute;
left:57px;
top:0px;
width:16px;
height:16px;
z-index:4;
background-color: #FF3300;
}
#apDiv69 {
position:absolute;
left:87px;
top:0px;
width:16px;
height:16px;
z-index:5;
}
#apDiv70 {
position:absolute;
left:117px;
top:0px;
width:16px;
height:16px;
z-index:6;
}
#apDiv71 {
position:absolute;
left:147px;
top:0px;
width:16px;
height:16px;
z-index:7;
}
#apDiv72 {
position:absolute;
left:180px;
top:3px;
width:13px;
height:12px;
z-index:8;
}
#apDiv73 {
position:absolute;
left:0px;
top:3px;
width:13px;
height:12;
z-index:9;
}

.ui-dialog
{
position:fixed;
}

-->
</style>
<script type="text/javascript">
<!--
function MM_findObj(n, d) { //v4.01
var p,i,x;  if(!d) d=document; if((p=n.indexOf("?"))>0&&parent.frames.length) {
d=parent.frames[n.substring(p+1)].document; n=n.substring(0,p);}
if(!(x=d[n])&&d.all) x=d.all[n]; for (i=0;!x&&i<d.forms.length;i++) x=d.forms[i][n];
for(i=0;!x&&d.layers&&i<d.layers.length;i++) x=MM_findObj(n,d.layers[i].document);
if(!x && d.getElementById) x=d.getElementById(n); return x;
}
function MM_preloadImages() { //v3.0
var d=document; if(d.images){ if(!d.MM_p) d.MM_p=new Array();
var i,j=d.MM_p.length,a=MM_preloadImages.arguments; for(i=0; i<a.length; i++)
if (a[i].indexOf("#")!=0){ d.MM_p[j]=new Image; d.MM_p[j++].src=a[i];}}
}
function MM_swapImgRestore() { //v3.0
var i,x,a=document.MM_sr; for(i=0;a&&i<a.length&&(x=a[i])&&x.oSrc;i++) x.src=x.oSrc;
}
function MM_swapImage() { //v3.0
var i,j=0,x,a=MM_swapImage.arguments; document.MM_sr=new Array; for(i=0;i<(a.length-2);i+=3)
if ((x=MM_findObj(a[i]))!=null){document.MM_sr[j++]=x; if(!x.oSrc) x.oSrc=x.src; x.src=a[i+2];}
}

$(document).ready(function()
{
if($.browser.mozilla == true)
{
if (screen.height<=1050)
{
$('.subitem-02').css('font-size','13px');
$('.titulo-oferta').css('height','30px');
}
}

$( "#catalogo" ).dialog({
autoOpen: false,
position: {at: "center top"},
width: 850,
height: 680
});

});
//-->
</script>
</head>
<body onload="MM_preloadImages('img/boton-webdesktop02.jpg','img/radio02.gif','img/fusion02.gif','img/tour02.gif','img/germina02.jpg','img/boton-acp02.jpg','img/boton-virtuales02.jpg')">
<div id="apDiv3">
<div id="apDiv18"></div>
<div id="apDiv4"><div id="apDiv8">
<div id="apDiv9">
<table width="135" border="0" cellspacing="0" cellpadding="4">
<tr>
<td><div align="center"><a href='https://www.facebook.com/ufgoficial' target='_blank'><img src="img/FB-logo.png" width="30" height="28" class='img-boton' /></a></div></td>
<td><div align="center"><a href='https://twitter.com/UFGOficial' target='_blank'><img src="img/twitter-logo.png" width="30" height="28"  class='img-boton' /></a></div></td>
<td><div align="center"><a href='http://www.youtube.com/user/redsocialufg?feature=mhw4' target='_blank'><img src="img/youtube-logo.png" width="30" height="28" class='img-boton' /></a></div></td>
<td><div align="center"><a href='http://punto105.com/' target='_blank'><img src="img/Link-Punto105-Radio.jpg" width="80" height="25" class='img-boton' /></a></div></td>
</tr>
</table>
</div>
<form id="fBusqueda" name="fBusqueda" style="padding:0px;margin:0px" action="buscador.php" method="post">
<div id="apDiv10">
<input id="txtBuscar" name="txtBuscar" style="width: 162px; height: 16px; background-color:e3e3e3; border: 1px solid #cccccc; font-size:10pt; color: #000000" type="text" value="">
</div>
<div id="apDiv11"><img src="img/boton-buscador.jpg" class="img-boton" height="20" width="25" onClick="document.getElementById('fBusqueda').submit()"></div>
</form>
<img src="img/logo-slogan.png" width="637" height="75" /></div>
<div class="help" id="apDiv12"><span onclick="openPopup('comentario','info.php?dst=1',400,350);">Información y contacto | Ayuda</span></div>
<div id="apDiv13"></div>
<div class="menu-arriba" id="apDiv14">
<table width="927" border="0" cellspacing="0" cellpadding="0">
<tr>
<td class="TD01" width="70" bgcolor="#FF6600"><div align="center" onClick="location.href='http://www.ufg.edu.sv/'">INICIO</div></td>
<td class="TD01" id="M,1" width="120"><div align="center" onClick="location.href='ini.nuestra.institucion.html'">NUESTRA INSTITUCIÓN</div></td>
<td class="TD01" id="M,2" width="119"><div align="center" onClick="location.href='ini.facultades.html'">FACULTADES</div></td>
<td class="TD01" id="M,3" width="135"><div align="center" onClick="location.href='ini.tecnologia.html'">TECNOLOGÍA</div></td>
<td class="TD01" id="M,4" width="137"><div align="center" onClick="location.href='ini.innovacion.html'">INNOVACIÓN</div></td>
<td class="TD01" id="M,5" width="121"><div align="center" onClick="location.href='ini.calidad.html'">CALIDAD</div></td>
<td class="TD01_1" id="M,6" width="225"><div align="center" onClick="location.href='http://comunidad.ufg.edu.sv/'">ACTIVIDAD ESTUDIANTIL</div></td>
</tr>
</table>
</div>
</div>
<div id="apDiv5"><div id="apDiv19">
<table width="191" border="0" align="center" cellpadding="0" cellspacing="0">
<tr>
<td height="36" class="titulo-oferta">Infórmate Ya</td>
</tr>
<tr>
<td height="10" class="TD03">[+] EGRESADOS Y GRADUADOS</td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://registro.ufg.edu.sv/InformacionEgresados/" class="subitem-02">» Curso básico para egresados</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://registro.ufg.edu.sv/InformacionEgresados/" class="subitem-02">» Especializaciones</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://registro.ufg.edu.sv/infografia_egreso/infografia_egreso.html" class="subitem-02" target="_blank">» Proceso de Graduación</a></td>
</tr>
<tr>
<td height="7"></td>
</tr>
<tr>
<td height="10" class="TD03">[+] POSTGRADOS UFG</td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://www.ufg.edu.sv/postgrados/palabras.html" class="subitem-02">» Maestrías</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://www.ufg.edu.sv/postgrados/palabras.html?1" class="subitem-02">» Solicitud de información</a></td>
</tr>
<tr>
<td height="7"></td>
</tr>
<tr>
<td height="10" class="TD03">[+] EDUCACIÓN CONTINUA</td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://www.ufg.edu.sv/ini.curdip.html?l=2&a=7&a=0&t=1" class="subitem-02">» Diplomados</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://www.ufg.edu.sv/ini.curdip.html?l=20&a=0&a=7&t=0" class="subitem-02">» Cursos</a></td>
</tr>
<tr>
<td height="7"></td>
</tr>
<tr>
<td height="10" class="TD03">[+] Servicios Universitarios</td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://www.ufg.edu.sv/su.ie.ayuwd.html" class="subitem-02">» Servicios Académicos</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="http://registro.ufg.edu.sv/carreras/asistencia_financiera" class="subitem-02">» Asistencia Financiera</a></td>
</tr>
<tr>
<td height="10" class="subitem-02"><a href="#" onClick="document.getElementById('fcatalogo').src='https://webdesktop.ufg.edu.sv/catalogo/index.html';$('#catalogo').dialog('open');" class="subitem-02">» Catálogo Institucional</a></td>
</tr>
</table>
</div>

<div id="apDiv20"><a href="https://webdesktop.ufg.edu.sv/" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image26','','img/BotonWebDesktop02.jpg',1)"><img src="img/BotonWebDesktop01.jpg" name="Image26" width="205" height="54" border="0" id="Image26" /></a></div>
<div id="apDiv57"><a href=" http://registro.ufg.edu.sv/carreras" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image24','','img/BotonCarreras.jpg',1)"><img src="img/BotonCarreras01.jpg" name="Image24" width="205" height="54" border="0" id="Image24" /></a></div>
<div id="apDiv21"><a href="http://registro.ufg.edu.sv/carrerasenlinea" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image20','','img/BotonEnLinea.jpg',1)"><img src="img/BotonEnLinea01.jpg" name="Image20" width="205" height="54" border="0" id="Image20" /></a></div>
<div id="apDiv62"><a href="http://biblioteca.ufg.edu.sv/" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image25','','img/BotonBibliotecario02.jpg',1)"><img src="img/BotonBibliotecario01.jpg" name="Image25" width="205" height="54" border="0" id="Image25" /></a></div>
<!--<div id="apDiv21"><a href="http://www.ufg.edu.sv/su.ie.ayuwd.html" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image24','','img/BotonUniversitarios02.jpg',1)"><img src="img/BotonUniversitarios01.jpg" name="Image24" width="205" height="54" border="0" id="Image24" /></a></div>-->
<div id="apDiv74"><a href="http://icti.ufg.edu.sv/" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image19','','img/BotonICTI02.jpg',1)"><img src="img/BotonICTI01.jpg" name="Image19" width="205" height="54" border="0" id="Image19" /></a></div>
<!--<div id="apDiv74"><a href="#" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image20','','img/btn_Catalogo2.jpg',1)"><img src="img/btn_Catalogo1.jpg" name="Image20" width="205" height="54" border="0" id="Image20" onClick="document.getElementById('fcatalogo').src='https://webdesktop.ufg.edu.sv/catalogo/index.html';$('#catalogo').dialog('open');" /></a></div>-->
<!--<div id="apDiv74"><a href="#" onmouseout="MM_swapImgRestore()" onmouseover="MM_swapImage('Image20','','img/boton_TVirtual02.jpg',1)"><img src="img/boton_TVirtual01.jpg" name="Image20" width="205" height="54" border="0" id="Image20" /></a></div>-->

<div id="apDiv22" class="texto-normal" style="position:absolute;">
<div class="titulo-encuesta"><img src="img/titulo_encuesta.fw.png" /></div>
<br>
<div id="cencuesta" style="margin:5px;text-align:justify">

<div style="margin:5px;text-align:justify">&iquest;Cree que la situaci&oacute;n del pa&iacute;s mejorar&aacute; con la realizaci&oacute;n de cambios en el Gabinete de Gobierno?</div><br>
<form class="formulario_encuesta" style="margin-top:0px;margin-bottom:0px" name="f_encuesta428" id="f_encuesta428" method="post" action="encuesta.php">
<input type="hidden" name="idencuesta" value="428"/>
<input type="hidden" name="tipo" value="R"/>
<input type="radio" name="op" value="1931">S&iacute;<br><input type="radio" name="op" value="1932">No<br><input type="radio" name="op" value="1933">A medias<br><input type="radio" name="op" value="1934">No sabe<br><input type="radio" name="op" value="1935">Le es indiferente<br><input name="ok" value="" type="submit" style="background-image:url('img/boton-votar.jpg');cursor:pointer;position:relative;left:68px;top:6px;width:46px;height:18px;border:0px;"><br><br></form>
</div>
</div>
</div>
<div id="apDiv6">
<div id="apDiv15"><img width="710" height="329" id="banner" />
<div id="apDiv31">
<div id="apDiv32" onclick="javascript:back_banner();"><img src="img/arrow-izq.gif" width="13" height="12" /></div>
<div class="div-numeros" id="cuadro-0" onclick="javascript:aqui_banner(0);">1</div>
<div class="div-numeros" id="cuadro-1" onclick="javascript:aqui_banner(1);">2</div>
<div class="div-numeros" id="cuadro-2" onclick="javascript:aqui_banner(2);">3</div>
<div class="div-numeros" id="cuadro-3" onclick="javascript:aqui_banner(3);">4</div>
<div class="div-numeros" id="cuadro-4" onclick="javascript:aqui_banner(4);">5</div>
<div class="div-numeros" id="cuadro-5" onclick="javascript:aqui_banner(5);">6</div>
<div id="apDiv38" onclick="javascript:next_banner();"><img src="img/arrow-der.gif" width="13" height="12" /></div>
</div>
<script language="javascript">
ini_banner('img/banner1.jpg||http://www.ufg.edu.sv/aniversario.html,img/banner2.jpg||http://www.ufg.edu.sv/aniversario.html,img/banner3.jpg||http://www.ufg.edu.sv/aniversario.html,img/banner4.jpg||http://www.ufg.edu.sv/aniversario.html,img/banner5.jpg||http://www.ufg.edu.sv/aniversario.html,img/banner6.jpg||http://www.ufg.edu.sv/aniversario.html');
</script>
</div>
<div id="apDiv16">
<br/>
<img src="img/barra_carteleraUFG.jpg"  />
</div>

<div id="apDiv28">
<div id="apDiv42"><img src="img/img_eventos.jpg"  /></div>
<div id="apDiv43"><img  width="400" height="245" id="news" /></div>
<div class="texto-normal" id="apDiv44">
</div>
<div id="apDiv45">
<div id="apDiv46"><img src="img/arrow-izq.gif" width="13" height="12" onclick="javascript:back_noticia();" /></div>
<div class="div-numeros2" id="cube-0" onclick="javascript:aqui_noticia(0);">1</div>
<div class="div-numeros2" id="cube-1" onclick="javascript:aqui_noticia(1);">2</div>
<div class="div-numeros2" id="cube-2" onclick="javascript:aqui_noticia(2);">3</div>
<div class="div-numeros2" id="cube-3" onclick="javascript:aqui_noticia(3);">4</div>
<div class="div-numeros2" id="cube-4" onclick="javascript:aqui_noticia(4);">5</div>
<div class="div-numeros2" id="cube-5" onclick="javascript:aqui_noticia(5);">6</div>
<div class="div-numeros2" id="cube-6" onclick="javascript:aqui_noticia(6);">7</div>
<div id="apDiv54"><img src="img/arrow-der.gif" width="13" height="12" onclick="javascript:next_noticia();" /></div>
</div>
<div class="texto-3noticias" id="apDiv55"></div>
<div class="mas-news" id="apDiv56"><a href="noticias.php?tipo=E">Más eventos [+]</a></div>
<script type="text/javascript">ini_noticia('img/c23db97965a87b3aa79f60678cfeac09.jpg||Vacaciones de Semana Santa 2018.||Ent&eacute;rate sobre las Vacaciones de Semana Santa 2018.||N.1352.html,img/5ab6a63ea026fc2da8954a572da89d3f.jpg||Diplomado en Administraci&oacute;n de la Cadena de Abastecimiento y Log&iacute;stica.||Inscr&iacute;base en el Diplomado en Administraci&oacute;n de la Cadena de Abastecimiento y Log&iacute;stica.||N.1331.html,img/f79c44aec60defced6552ba0941a2c8e.jpg||Curso de Auditores Internos en Sistema de Calidad ISO 9001:2015.||Inscr&iacute;bete Curso de Auditores Internos en Sistema de Calidad ISO 9001:2015||N.1334.html,img/6feef3daccdede6caac8fbbd6fa04282.jpg||Descubre tu pasi&oacute;n con la UFG.||Descubre tu pasi&oacute;n con la UFG - Proceso de Orientaci&oacute;n Vocacional.||N.1291.html,img/76316e805d540b69bdc82e12d8efcc3d.jpg||Solemnes Actos de Graduaci&oacute;n UFG 2018.||Ent&eacute;rate sobre Los Solemnes Actos de Graduaci&oacute;n UFG 2018.||N.1281.html,img/7baaa887f8ea256eb970949c62a28e9e.jpg||Prevengamos la Conjuntivitis||Prevengamos la Conjuntivitis||N.1192.html,img/386a4ebd4057cadfdff6c7b86e6bc343.jpg||Tarjeta Estudio Prom&eacute;rica||Tarjeta Estudio Prom&eacute;rica. Solic&iacute;tala.||N.1219.html||')</script>
</div>

<div id="apDiv29">
<div id="apDiv39"><img src="img/img_noticias.jpg"/></div>
<div id="apDiv40">
<table width="240" border="0" cellspacing="3" cellpadding="2">
<tr id="tr1"></tr>
<tr id="tr2"></tr>
<tr id="tr3"></tr>
<tr id="tr4"></tr>
<tr id="tr5"></tr>
<tr id="tr6"></tr>
<tr id="tr7"></tr>
<tr id="tr8"></tr>
<tr id="tr9"></tr>
<tr id="tr10"></tr>
<tr id="tr11"></tr>
<tr id="tr12"></tr>
<tr id="tr13"></tr>
<tr id="tr14"></tr>
<tr id="tr15"></tr>
</table>
</div>
<div class="mas-news" id="apDiv41"><a href="noticias.php?tipo=N">Más noticias [+]</a></div>
<script type="text/javascript">ini_evento('4 Dic.||Concurso de Oratoria en Ingl&eacute;s||E.1270.html;;15 Nov.||Semana de la Salud Mental.||E.1234.html;;14 Nov.||Ganador de TV 32" en Tabling UFG.||E.1235.html;;19 Oct.||Beneficios UFG con Grupo Premium.||E.1184.html;;19 Oct.||Ganador en Tabling UFG Credomatic||E.1181.html;;13 Ene.||I Promoci&oacute;n UFG 2016||E.919.html;;13 Ene.||II Promoci&oacute;n UFG 2016||E.921.html;;13 Ene.||III Promoci&oacute;n UFG 2016||E.923.html;;13 Ene.||IV Promoci&oacute;n UFG 2016||E.924.html;;28 Oct.||Ganadoras del V Concurso de Oratoria en Idioma Ingl&eacute;s||E.856.html;;20 Oct.||XXVI edici&oacute;n del Foro Aportando Soluciones: "An&aacute;lisis de la competitividad y desarrollo econ&oacute;mico de El Salvador".||E.847.html;;26 Sep.||III Seminario: "Caracter&iacute;sticas y medidas de seguridad de los d&oacute;lares y funciones de un cajero de banco"||E.829.html;;21 Sep.||"Salarru&eacute; en el per&iacute;odo Patria".||E.826.html;;6 Jul.||D&iacute;a del Maestro UFG 2016||E.770.html;;3 Jun.||V Concurso de Litigaci&oacute;n Oral||E.744.html;;5 May.||Estudiantes UFG representan a El Salvador.||E.677.html;;30 Abr.||V&iacute;ctima del phubbing||E.623.html;;30 Abr.||Regal&iacute;as por Derechos de Autor.||E.622.html;;25 Feb.||UFG inaugura su Centro de Modelaje Matem&aacute;tico ?Carlos Castillo-Ch&aacute;vez?||E.613.html;;19 Feb.||Crezcamos para unirnos||E.608.html;;19 Feb.||La Verdad...||E.607.html;;10 Feb.||Concurso InterUniversitario de Dise&ntilde;o de Edificio Ecol&oacute;gico||E.603.html;;9 Feb.||Presentaci&oacute;n del libro "El Refuerzo Educativo"||E.601.html;;8 Feb.||VII Entrega Anual de Becas Universitarias||E.592.html;;12 Ene.||Un modelo &oacute;ptimo en la Educaci&oacute;n salvadore&ntilde;a||E.584.html;;9 Ene.||Celebraciones Navide&ntilde;as UFG 2015.||E.583.html;;8 Ene.||La Lectura: mi compromiso de 2016.||E.581.html;;15 Dic.|| XIII Concurso Interuniversitario sobre Competencias para Juicios Orales en Justicia Penal Juvenil - 2015||E.576.html;;19 Oct.||Rally Latinoamericano de Innovaci&oacute;n||E.538.html;;7 Oct.||Escribir bien ¿para qu&eacute;?: La necesidad de una comunicaci&oacute;n efectiva a trav&eacute;s del discurso escrito.||E.532.html;;18 Sep.||Bases del Concurso de Ideas y Modelos de Negocios para Estudiantes UFG.||E.491.html;;31 Ago.||M&aacute;s Cub&iacute;culos de Estudio Grupal en las Bibliotecas UFG||E.497.html;;26 Jun.||Foro Internacional contra la Violencia Escolar||E.472.html;;4 Jun.||Libro: Democracia y Financiamiento de Partidos Pol&iacute;ticos||E.471.html;;3 Jun.||Ganadores del IV Concurso de Litigaci&oacute;n Oral.||E.469.html;;30 Abr.||Acceso Peatonal habilitado entre la Avenida Ol&iacute;mpica y la 57 Av. Sur||E.379.html;;28 Abr.||Selecci&oacute;n de F&uacute;tbol Playa UFG||E.424.html;;15 Abr.||Conferencia "La Historia del Internet en El Salvador"||E.413.html;;31 Ene.||Lanzamiento UFG Online University||E.292.html;;21 Ene.||Entrega de Becas UFG BAC Credomatic 2015||E.350.html;;15 Ene.||Firma de Carta de Entendimiento UFG - Entrepreneurs Organization Cap&iacute;tulo El Salvador||E.346.html;;16 Dic.||Felicitaci&oacute;n por Investidura Acad&eacute;mica Doctoral||E.331.html||')</script>
</div>
<div id="apDiv30"><img src="img/division.jpg" width="1" height="240" /></div>
</div>
<div id="apDiv7">
<div align="center">
<table width="927" border="0" cellspacing="0" cellpadding="0">
<tr>
<td width="463" height="95"><img src="img/pie-pagina.jpg" width="463" height="95" /></td>
<td width="464" height="95" class="texto-piepagina">
<p>Nuevo Ingreso San Salvador | Edificio de Atención al Estudiante,<br/>1er. Nivel, Condominio Centro Roosevelt, 55 Av. Sur,<br/>Entre Alameda Roosevelt y Av. Olímpica. Tel. 2209-2816, 2209-2839</p>
<p>Copyright © 2014 UFG | Calle El Progreso No. 2748, Edificio de Rectoría<br>San Salvador, El Salvador. Tel. 2249-2700</p>
<p>Centro Regional de Occidente | Final 9a. Calle Poniente, entre 18 y 20 <br>Av. Sur, Santa Ana. Tel. 2441-2927, 2447-3403</p>
</td>
</tr>
</table>
</div>
<map name="calidad">
<area shape=rect coords="4,4,87,85" href="http://www.mined.gob.sv/cda/convocatorias.htm" target="_blank">
<area shape=rect coords="96,20,130,74" href="http://www.ufg.edu.sv/lsqa.html" target="_blank">
<!--<area shape=rect coords="110,10,214,54" href="http://www.ufg.edu.sv/Qualityaustria.html" target="_blank">
<area shape=rect coords="216,0,269,56" href="http://www.ufg.edu.sv/Qualityaustria.html" target="_blank">-->
</map>
</div>
<div id="apDiv61"></div>

<div id="apDiv78">
<div id="apDiv79">
<div id="apDiv80"><img src="img/loguito-UFG.jpg" width="54" height="19" /></div>
</div>
<div class="interlineado-texto" id="apDiv82">
<table width="150" border="0" cellspacing="0" cellpadding="0">
<tr>
<td height="18" class="texto-celeste">Nuestra instituci&oacute;n</td>
</tr>

<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/nuestra.historia.html">Nuestra historia</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/mision.vision.valores.html">Misi&oacute;n, visi&oacute;n y valores</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/politicas.de.calidad.html">Pol&iacute;ticas de calidad</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/rectoria.html">Mensaje del Rector</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/c.acdayacaai.html">Acreditaciones de calidad</a></td>
</tr>
<!-- <tr>
<td class="texto-mapa"><a href="" >Plan estrat&eacute;gico UFG</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="" >Normas y reglamentos</a></td>
</tr> -->
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/catalogo-ufg.html" >Cat&aacute;logo institucional</a></td>
</tr>

<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/est.org.html">Estructura organizacional</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/convenios.html">Convenios</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/evolydes.html">Evoluci&oacute;n y desarrollo</a></td>
</tr>
</table>
</div>
<div id="apDiv83">
<table width="165" border="0" cellspacing="0" cellpadding="0">

<tr>
<td class="texto-mapa"><span class="texto-celeste">Facultades</span></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://fad.ufg.edu.sv/">Arte y Dise&ntilde;o</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://fce.ufg.edu.sv/">Ciencias Econ&oacute;micas</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://fcj.ufg.edu.sv/">Ciencias Jur&iacute;dicas</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://fcs.ufg.edu.sv/">Ciencias Sociales</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://fis.ufg.edu.sv/">Ingenier&iacute;a y Sistemas</a></td>
</tr>

<tr>
<td height="15" class="texto-mapa"></td>
</tr>
<tr>
<td height="10" class="texto-normal"><span class="texto-celeste">Tecnolog&iacute;a</span></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/inftecn.html">Infraestructura tecnol&oacute;gica</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/lab.html">Laboratorios</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/serelin.html">Servicios en l&iacute;nea</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/teceduc.html">Tecnolog&iacute;a educativa</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/acadtec.html">Academias de tecnolog&iacute;a</a></td>
</tr>
</table>
</div>
<div id="apDiv84">
<table width="170" border="0" cellpadding="0" cellspacing="0" class="texto-normal">
<tr>
<td class="texto-celeste">Actividad estudiantil</td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://comunidad.ufg.edu.sv/becas.html" >Becas</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://comunidad.ufg.edu.sv/deporte.html">Deportes</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://comunidad.ufg.edu.sv/extension.cultural.html">Extensi&oacute;n cultural</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://comunidad.ufg.edu.sv/orientacion.vocacional.html">Orientaci&oacute;n vocacional</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://comunidad.ufg.edu.sv/servicio.social.estudiantil.html">Servicio social estudiantil</a></td>
</tr>
<tr>
<td height="15" class="texto-normal">&nbsp;</td>
</tr>
<tr>
<td class="texto-mapa"><span class="texto-celeste">Otros enlaces</span></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.universia.com.sv/">Universia</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://telescopi.upc.edu/">Telescopi</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.raices.org.sv/">Raices</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.tecoloco.com.sv/">Tecoloco</a></td>
</tr>
<!-- <tr>
<td class="texto-mapa"><a href="http://www.gradodigital.edu.sv/">Grado Digital</a></td>
</tr> -->
</table>
</div>
<div id="apDiv85">
<table width="165" border="0" cellspacing="0" cellpadding="0">
<tr>
<td height="10" class="texto-mapa"><span class="texto-celeste">Innovaci&oacute;n</span></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/i.vinuivemp.html">Relaci&oacute;n Universidad-Empresa</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/i.germina.html">Incubadora  GERMINA</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/i.cdmype.ufg.html">CDMYPE-UFG</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/i.icti.ufg.html">ICTI</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/i.proysoc.html">Proyecci&oacute;n social</a></td>
</tr>
<tr>
<td height="15" class="texto-mapa"></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><span class="texto-celeste">Calidad</span></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><span class="texto-mapa"><a href="http://www.ufg.edu.sv/c.acdayacaai.html">Acreditaciones: CdA y ACAAI</a></span></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><span class="texto-normal"><a href="http://www.ufg.edu.sv/c.niso.html">Norma ISO 9001:2008</a></span></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/c.ayrufg.html">Asociaciones y redes a las que pertenece la UFG</a></td>
</tr>
<tr>
<td height="10" class="texto-mapa"><a href="http://www.ufg.edu.sv/c.pacp.html">Programa ACP</a></td>
</tr>
</table>
</div>
<div id="apDiv86">
<table width="130" border="0" cellspacing="0" cellpadding="0">
<tr>
<td class="texto-celeste">Nuestras carreras</td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://nuevoingreso.ufg.edu.sv" >Carreras</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://nuevoingreso.ufg.edu.sv/ni.requisitos.html">Requisitos</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://nuevoingreso.ufg.edu.sv/ni.aranceles.html">Aranceles</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://nuevoingreso.ufg.edu.sv/ni.calendario.html">Calendarios y horarios</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://registro.ufg.edu.sv/InformacionEgresados/">Curso para egresados</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://registro.ufg.edu.sv/InformacionEgresados/">Especializaciones</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/postgrados/palabras.html">Maestr&iacute;as</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://www.ufg.edu.sv/postgrados/palabras.html" >Informaci&oacute;n maestr&iacute;as</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://diplomados.ufg.edu.sv/">Diplomados</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://cursos.ufg.edu.sv/">Cursos</a></td>
</tr>
<tr>
<td class="texto-mapa"><a href="http://seminarios.ufg.edu.sv/">Seminarios</a></td>
</tr>
</table>
</div>
</div>
</div>
</div>

<div id="catalogo" title="Catálogo Institucional UFG">
<iframe id="fcatalogo" width="100%" height="670" frameborder="no" src="" style="border: 0px solid black;"></iframe>
</div>


<!-- Piwik -->
<script type="text/javascript">
var _paq = _paq || [];
_paq.push(["trackPageView"]);
_paq.push(["enableLinkTracking"]);

(function() {
var u=(("https:" == document.location.protocol) ? "https" : "http") + "://analytics.ufg.edu.sv/";
_paq.push(["setTrackerUrl", u+"piwik.php"]);
_paq.push(["setSiteId", "2"]);
var d=document, g=d.createElement("script"), s=d.getElementsByTagName("script")[0]; g.type="text/javascript";
g.defer=true; g.async=true; g.src=u+"piwik.js"; s.parentNode.insertBefore(g,s);
})();
</script>
<!-- End Piwik Code -->

</body>
</html>