

<!DOCTYPE html>
<html>
<head>
    <script type="text/javascript" src="/ruxitagentjs_ICA2SVfqr_10139180201161915.js" data-dtconfig="rid=RID_2418|rpid=1801393093|domain=tecoloco.com.sv|reportUrl=/rb_bf05879vqo|featureHash=ICA2SVfqr|lastModification=1521316405617|dtVersion=10139180201161915|tp=500,50,0,1|agentUri=/ruxitagentjs_ICA2SVfqr_10139180201161915.js"></script><link href='https://fonts.googleapis.com/css?family=Open+Sans:400,300,600' rel='stylesheet' type='text/css'>
    <link href="/Content/2016/font-awesome.min.css" rel="stylesheet"/>

    <meta charset="utf-8">
    <!-- IE Edge Meta Tag -->
    <meta http-equiv="X-UA-Compatible" content="IE=edge"> 




    <meta name="viewport" content="width=device-width, initial-scale=1, user-scalable=no">

    <link rel="icon" href="/Content/images/favicon.ico" type="image/x-icon" />
    
    <title>Trabajo en El Salvador Empleo en El Salvador www.tecoloco.com.sv</title>
    

    

    <script src="/Scripts/2016/modernizr-2.6.2.js"></script>
    <script src="/Scripts/PLNativeBridge_v2.js"></script>


    <link rel="stylesheet"  href="/Content/themes/base/jquery-ui.css" type="text/css" />    
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/bootstrap.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/bootstrap-responsive.css" type="text/css" />

    <link rel="stylesheet" media='screen and (max-width: 1023px)' href="https://maxcdn.bootstrapcdn.com/bootstrap/3.3.5/css/bootstrap.min.css">
    <link rel="stylesheet" media='screen and (max-width: 1023px)' href="/Content/2016/responsive2016/responsive.css">
    <link rel="stylesheet" media='screen and (max-width: 1023px)' href="/Content/2016/responsive2016/default-color.css">
    <link rel="stylesheet" media='screen and (max-width: 1023px)' href="/Content/2016/responsive2016/reset-old-style.css">

    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/tecoloco.css?v=2.25" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/themes/base/jquery.ui.datepicker.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/Site.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/styles.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/kendo/kendo.common.min.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/kendo/kendo.default.min.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/kendo/kendo.silver.min.css" type="text/css" />
    <link rel="stylesheet" media='screen and (min-width: 1024px)' href="/Content/estilosprite.css" type="text/css" />

    




    <!-- Optional IE8 Support -->
    <!--[if lt IE 9]>
      <script src="https://oss.maxcdn.com/html5shiv/3.7.2/html5shiv.min.js"></script>
      <script src="https://oss.maxcdn.com/respond/1.4.2/respond.min.js"></script>
    <![endif]-->
    

    <!-- jQuery -->
    <script src="https://ajax.googleapis.com/ajax/libs/jquery/1.11.3/jquery.min.js"></script>
    <script src="https://code.jquery.com/jquery-migrate-1.4.0.js"></script>
    <script src="/Scripts/2016/responsive/responsive.js"></script>



    <!-- Minified JavaScript -->
    <script src="https://maxcdn.bootstrapcdn.com/bootstrap/3.3.5/js/bootstrap.min.js"  ></script>

          
          




    


    
    
    <script src="/Scripts/jquery-ui-dev/jquery.ui.core.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.datepicker.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.widget.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.button.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.dialog.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.mouse.js"></script>

    <script src="/Scripts/jquery-ui-dev/jquery.ui.draggable.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.position.js"></script>
    <script src="/Scripts/jquery-ui-dev/jquery.ui.resizable.js"></script>
    <script src="/Scripts/jquery.ui.datepicker-es.js"></script>



    <script src="/Scripts/jquery.validate.js"></script>
    <script src="/Scripts/jquery.validate.unobtrusive.js"></script>


    <script src="/Scripts/knockout-2.1.0.js"></script>
    
    <script src="/Scripts/knockout.validation.js"></script>


    
    <script src="/Scripts/moment.js"></script>
    <script src="/Scripts/jquery.blockUI.js"></script>
    <script src="/Scripts/jquery.cookie.js"></script>

    
    <script src="/Scripts/kendo/custom/kendo.core.js"></script>
    <script src="/Scripts/kendo/custom/kendo.fx.js"></script>
    <script src="/Scripts/kendo/custom/kendo.userevents.js"></script>
    <script src="/Scripts/kendo/custom/kendo.draganddrop.js"></script>
    <script src="/Scripts/kendo/custom/kendo.window.js"></script>

    <script src="/Scripts/TecolocoScripts.js"></script>
    <script src="/Scripts/tecoloco.js"></script>
    <script src="/Scripts/navCvs.js"></script>
    <script src="/Scripts/jquery.pngFix.js"></script>
    <script src="/Scripts/bpopup.js"></script>    


    <script src="/Scripts/knockout.mapping-latest.debug.js"></script>






          
            <link rel="alternate" href="android-app://com.stepstone.tecoloco/sttl/source/homepage" />
        






    <!-- Google Analityc -->
    <script type="text/javascript">
        //<![CDATA[
        var gaJsHost = (("https:" == document.location.protocol) ? "https://ssl." : "http://www.");
        document.write(unescape("%3Cscript src='" + gaJsHost + "google-analytics.com/ga.js' type='text/javascript'%3E%3C/script%3E"));
        //]]>
    </script>
    <script type="text/javascript">
        //<![CDATA[
        try {
            var pageTracker = _gat._getTracker('UA-2829140-17');
            pageTracker._trackPageview();
        } catch (err) { }
        //]]>
    </script>
    
    <!-- Google Tag Manager -->
    <script>(function(w,d,s,l,i){w[l]=w[l]||[];w[l].push({'gtm.start':
            new Date().getTime(),event:'gtm.js'});var f=d.getElementsByTagName(s)[0],
            j=d.createElement(s),dl=l!='dataLayer'?'&l='+l:'';j.async=true;j.src=
            'https://www.googletagmanager.com/gtm.js?id='+i+dl;f.parentNode.insertBefore(j,f);
    })(window,document,'script','dataLayer','GTM-NCMWQ3X');</script>
    <!-- End Google Tag Manager -->


    

    <style>

        #fade { 
  /* Blacks out content during ad display. A hat tip to Brett DeWoody of Digital Wax Works (http://www.DigitalWaxWorks.com) for this piece... */
  display: none;
  background-color: #000;
  position: fixed; 
  left: 0; 
  top: 0;
  width: 100%; height: 100%;
  opacity: .70;
  z-index: 1000000;
}

#popupBlock {/* Sets positioning for ad... */
  display: none;
  float: left;
  position: fixed;
  top: 0; 
  left: 0;
  z-index: 1000001;
}

.sponsorad { /*These properties make the interstitial ad responsive*/
  border: 3px solid white;
  background: url('../img/red800.png');
  background-size: 90% auto;
  background-repeat: no-repeat;
  background-position: center 40%;
  padding: 3px; 
  position: fixed;
  top: 7.5%;
  left: 7.5%;
  width: 85%;
  height: auto;
  min-height: 85%;
  background-color: #CFCFCF;
  color: #5E5E5E
}


.sponsorad span { /*Styling for the phrase "A message from this week's sponsor..." */
  position: absolute;
  top: 1em;
  left: 1em;
  font-style: italic;
  max-width: 60%;
}

.sponsorad a:link { /* Styling the "close" link... */
  color: #5E5E5E;
  position: absolute;
  top: 1em;
  right: 1em;
  margin-left: 3em;
}

    </style>




</head>

    <body class=" " >
    <!-- Google Tag Manager (noscript) -->
    <noscript><iframe src="https://www.googletagmanager.com/ns.html?id=GTM-NCMWQ3X"
                      height="0" width="0" style="display:none;visibility:hidden"></iframe></noscript>
    <!-- End Google Tag Manager (noscript) -->
        <div class="visible-phone">


            <span class="clear"></span>
        </div>

        <div class="" >





            <noscript>
    <div class="jswarningdisabledontop">
        Para poder tener una mejor experiencia en la navegabilidad de nuestro sitio es necesario que habilites el uso de javascript en tu navegador.<br />  Para averiguar si el explorador admite JavaScript o para permitir las secuencias de comandos, consulte la ayuda en pantalla del explorador.
    </div>
</noscript>




            <div class="visible-phone mobile-menu ">
                <div class="mobile-main-menu-bar">
                    <a class="phone-btnBack btn-menu" onclick="goBack()">
                    </a>
                   
                    <a class="logo21" href="/">
                        
                    </a>
                    <a class="phone-btnMenuAux btn-menu itemT" data-toggle="collapse" data-target="#menuPrincipal"></a>
                    <span class="clear"></span>
                </div>


                <div id="menuPrincipal" class="collapse mobile-sub-menu">



                    <a class="phone-menu-item" href="/Default2.aspx"><span class="phone-icoTrabajos btn-menu"></span>Trabajos</a>
                    <a class="phone-menu-item" href="/contacto.aspx    "><span class="phone-icoContactos btn-menu"></span>Contactos</a>



                        <a class="phone-menu-item" href="/listado/empresas-destacadas.aspx"><span class="phone-icoStands btn-menu"></span>Empresas</a>
                    <a class="phone-menu-item" href="/blog"><span class="phone-icoBlog btn-menu"></span>Blog</a>



                        <a class="phone-menu-item" href="/frmQSomos.aspx"><span class="phone-icoInterrogante btn-menu"></span>Nosotros</a>




                        <a class="phone-menu-item" href="/empresas/testimoniales-de-empresas"><span class="phone-icoComillas btn-menu"></span>Testimonios</a>



                        <a class="phone-menu-item" href="/frmPreguntas.aspx"><span class="phone-icoAyuda1 btn-menu"></span>Preguntas</a>


                        <a href="/frmFeed.aspx" class="phone-menu-item"><span class="phone-icoRss btn-menu"></span>RSS Feed</a>



                    



                    <span class="clear"></span>
                </div>







                <span class="clear"></span>


                    <div class="mobile-main-menu-bar">

                        
    <a class="phone-btnSearch-sub2 btn-menu-sub1"></a>


                        <a class="phone-btnUser-sub1 btn-menu-sub1 itemT" data-toggle="collapse" data-target="#menuUsuario"></a>
                        <span class="clear"></span>
                    </div>
                    <div id="menuUsuario" class="collapse mobile-sub-menu">




                        <a class="phone-menu-item" href="/Candidate"><span class="phone-icoConfiguracion btn-menu"></span>Mi Cuenta</a>



                            <a id="IniciarSesion_HR" class="phone-menu-item" href="/Candidatos/frmAbreCuenta.aspx" target="_self"><span class="phone-icoNuevoUsuario btn-menu"></span>Reg&iacute;strate</a>


                        




                        <a class="phone-menu-item" href="javascript:getFeedData();"><span class="phone-icoSugerencias btn-menu"></span>Sugerencias</a>


                        <a class="phone-menu-item"><span class="phone-icoVacio btn-menu"></span></a>




                        <span class="clear"></span>
                    </div>
            </div>

            <span class="clear"></span>
            <br />



            <span class="clear"></span>


            <span class="clear"></span>
            <div class="container-fluid">
                <div class="header row-fluid hidden-phone">
                    <div class="pull-left">
                        <a class="logoTecoloco" href="/">
                            <img id="imgLogo" title="encuentra trabajos empleos vacantes y oportunidades laborales" class="logo" src="/Content/logos/tecoloco-ElSalvador.png" style="border-width: 0px;" />
                        </a>

                                    <h1>TRABAJOS EN EL SALVADOR Y EMPLEOS EN EL SALVADOR CON WWW.TECOLOCO.COM.SV</h1>
                                    <p>Encuentra las mejores ofertas de trabajo y ofertas de empleo en El Salvador con www.tecoloco.com.sv.</p>

                    </div>


    
    <a class="enlace" target="_blank"  href='/Home/SetClickAds?idAds=6sWJmYqnDsg%253d'>
                                            <img class="enlace" src="//content.tecoloco.com/Assets/publicidad/lxxpwlcp.5btDIGICEL_AD.jpg" style="border: 0">
                                        </a>

                </div>


                <nav class="row-fluid hidden-phone">
                    <div class="span12 menu">
                            <div id="comenzar">
                                <ul>
                                    <li>
<span class="sprite-btnLoginUser-align sprite-btnLoginUser"><a id="IniciarSesion_HI" href="/login.aspx">Inicio Candidatos</a></span>
                                        
                                    </li>

                                    <li class="visible-desktop">
                                            <a id="IniciarSesion_HR" href="/Candidatos/frmAbreCuenta.aspx" target="_self" class="sprite-btnRegistroUser-align sprite-btnRegistroUser">Regístrate</a>
                                    </li>

                                </ul>
                            </div>
<ul class="main"><li class="sprite-btnInicio"><a href="/">Inicio</a></li>
           <li class="sprite-btnTrabajos"><a id="hlBusqueda" href="/Default2.aspx">Trabajos</a></li> 
            <li class="visible-desktop sprite-btnBlog" id="btnBlog"><a id="hlBlog" title="Blog" href="/blog" target="_blank">Blog</a></li> 
   
<li class="sprite-btnContacto"><a id="hlContactos" href="/contacto.aspx">Contactos</a></li>    
    <li class="empresas-tecoloco visible-desktop btnEmpresas-align sprite-btnEmpresas"><a id="hlEmpresas" href="/loginEmpresas.aspx" target="_blank">Acceso<br />Empresas</a></li>
    
</ul>

                    </div>

                </nav>




                <nav class="row-fluid hidden-phone">

                    <ul class="sitemap span12">
                        <li class="ico sprite-icoSiteMap"></li>
                                <li>
                                    <a><div style='height: 20px;' class='svF'></div></a>
                                </li>
                                <li class="separador"></li>
                                <li>
                                    <a href="https://www.tecoloco.com.sv">www.tecoloco.com.sv</a>
                                </li>
                                <li class="separador"></li>
                    </ul>
                </nav>

                <div class="contenido-principal">



                    <div class="sidebar visible-desktop">
                        


<!--div class="titulo-landing"-->
<div class="imgTitLanding-align sprite-imgTitLanding">
    búsqueda por área
</div>
<div class="contenido-landing">
                <a href="/empleo-marketing-ventas">Mercadeo | Ventas (280)</a>
                <a href="/empleo-contabilidad">Finanzas | Contabilidad | Auditor&#237;a (160)</a>
                <a href="/empleo-informatica-internet">Inform&#225;tica | Internet (113)</a>
                <a href="/empleo-banco-servicios-financieros">Banca | Servicios Financieros (87)</a>
                <a href="/empleo-ingenieria-calidad">Producci&#243;n | Ingenier&#237;a | Calidad (86)</a>
                <a href="/empleo-restaurantes">Restaurantes (84)</a>
                <a href="/empleo-cualquier-area">Cualquier &#193;rea (69)</a>
                <a href="/empleo-mantenimiento">Mantenimiento (57)</a>
                <a href="/empleo-administrativo">Administraci&#243;n (48)</a>
                <a href="/empleo-oficinas">Apoyo de Oficina (48)</a>
                <a href="/empleo-profesionales">Puestos Profesionales (47)</a>
                <a href="/empleo-otros-trabajos">Varios (45)</a>
                <a href="/empleo-logistica">Operaciones | Log&#237;stica (42)</a>
                <a href="/empleo-recursos-humanos">Recursos Humanos (35)</a>
                <a href="/empleo-publicidad">Publicidad | Comunicaciones | Servicios (34)</a>
                <a href="/empleo-call-center">Call Center (29)</a>
                <a href="/empleo-bodega-almacenamiento">Almacenamiento (24)</a>
                <a href="/empleo-compras">Compras (21)</a>
                <a href="/empleo-salud">Salud (19)</a>
                <a href="/empleo-telefonia-telecomunicaciones">Telecomunicaciones (5)</a>

    <span class="clear"></span>
</div>

    <div class="foo-landing">
</div>
    <!--div class="titulo-landing"-->
    <div class="imgTitLanding-align sprite-imgTitLanding">
        búsqueda por cargo
    </div>
    <div class="contenido-landing">
                <a href="/empleo/ejecutivo-de-ventas">Ejecutiv@ de Ventas (72) </a>
                <a href="/empleo/cualquier-cargo">Cualquier Cargo (69) </a>
                <a href="/empleo/analista-programador">Analista | Programador (58) </a>
                <a href="/empleo/asistente-contable">Asistente Contable (39) </a>
                <a href="/empleo/chofer">Chofer (28) </a>
                <a href="/empleo/gestor-de-cobros">Gestor de Cobros (26) </a>
                <a href="/empleo/vendedor-rutero">Vendedor Rutero (25) </a>
                <a href="/empleo/cocinero">Cocinero (24) </a>
                <a href="/empleo/vendedor">Vendedor (23) </a>
                <a href="/empleo/analista-de-sistemas">Analista de Sistemas (18) </a>
                <a href="/empleo/repartidor">Repartidor (18) </a>
                <a href="/empleo/supervisor-de-produccion">Supervisor de Producci&#243;n (18) </a>
                <a href="/empleo/supervisor-de-ventas">Supervisor de Ventas (18) </a>
                <a href="/empleo/gerente-de-restaurante">Gerente de Restaurante (17) </a>
                <a href="/empleo/cajero">Cajer@ (14) </a>
                <a href="/empleo/ejecutivo-de-cuenta">Ejecutiv@ de Cuenta (14) </a>
                <a href="/empleo/mensajero">Mensajero (14) </a>
                <a href="/empleo/administrador">Administrador (13) </a>
                <a href="/empleo/asistente-administrativo">Asistente Administrativo (13) </a>
                <a href="/empleo/ejecutivo-pyme">Ejecutiv@ Pyme (13) </a>
                <a href="/empleo/jefe-de-sucursal-agencia">Jefe de Sucursal | Agencia (13) </a>
                <a href="/empleo/ejecutivo-de-banco">Otros Puestos Bancarios (13) </a>
                <a href="/empleo/asistente-de-recursos-humanos">Asistente de Recursos Humanos (12) </a>
                <a href="/empleo/contador-general">Contador General (12) </a>
                <a href="/empleo/ejecutivo-de-servicio-al-cliente">Ejecutiv@ de Servicio al Cliente (12) </a>
        <span class="clear"></span>
    </div>

<div class="foo-landing">
</div>
<!--div class="titulo-landing"-->
<div class="imgTitLanding-align sprite-imgTitLanding">
        <label>búsqueda por rubro</label> 
</div>
<div class="contenido-landing">
                <a href="/trabajo-servicios">Servicios (295) </a>
                <a href="/trabajo-comercial">Comercial (163) </a>
                <a href="/trabajo-bancos-financieras">Bancos | Financieras (147) </a>
                <a href="/trabajo-industrial">Industrial (143) </a>
                <a href="/trabajo-hoteleria-turismo-restaurantes">Hoteler&#237;a | Turismo | Restaurantes (88) </a>
                <a href="/trabajo-consumo-masivo-bebidas-alimentos-etc">Consumo Masivo (Bebidas | Alimentos) (55) </a>
                <a href="/trabajo-publicidad-marketing-rrpp">Publicidad | Marketing | RRPP (47) </a>
                <a href="/trabajo-agencia-de-reclutamiento">Agencia de Reclutamiento (45) </a>
                <a href="/trabajo-comercio-mayorista-intermediac-dist">Comercio Mayorista (Intermediac. | Dist.) (42) </a>
                <a href="/trabajo-logistica-distribucion">Log&#237;stica | Distribuci&#243;n (36) </a>
                <a href="/trabajo-consultoria-asesoria">Consultor&#237;a | Asesor&#237;a (35) </a>
                <a href="/trabajo-servicios-financieros-varios">Servicios Financieros Varios (25) </a>
                <a href="/trabajo-telecomunicaciones">Telecomunicaciones (24) </a>
                <a href="/trabajo-tecnologias-de-informacion">Tecnolog&#237;as de Informaci&#243;n (22) </a>
                <a href="/trabajo-servicios-varios">Servicios Varios (21) </a>
    
    <span class="clear"></span>
</div>
<div class="foo-landing">
</div>
                                <br /><h2 class="EmpresasReclutantesTit">Empresas que reclutan con nosotros:</h2>
                                <div id="empresas-destacadas">
                                    

                                    
<div id="content-empresas-destacadas">
    
<span>
                <a id="StandsControl1_d_ct100_h" href="/empresas-destacadas/trabajos-en-global-outsourcing_1633.aspx" >
                    <img id="StandsControl1_d_ct100_Image1" src="/stands.axd?image=GLobal-outsorcing-sv.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct101_h" href="/empresas-destacadas/trabajos-en-pollo-campero_515.aspx" >
                    <img id="StandsControl1_d_ct101_Image1" src="/stands.axd?image=logo-nuevo-pollo-camperooo.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct102_h" href="/empresas-destacadas/trabajos-en-almacenes-siman_512.aspx" >
                    <img id="StandsControl1_d_ct102_Image1" src="/stands.axd?image=nq4wghfh.vn0Siman-principal.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct103_h" href="/empresas-destacadas/trabajos-en-contactos-y-oportunidades_1309.aspx" >
                    <img id="StandsControl1_d_ct103_Image1" src="/stands.axd?image=contact stand.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct104_h" href="/empresas-destacadas/trabajos-en-forza-sa-de-cv_1303.aspx" >
                    <img id="StandsControl1_d_ct104_Image1" src="/stands.axd?image=forza stand.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct105_h" href="/empresas-destacadas/trabajos-en-banco-davivienda_502.aspx" >
                    <img id="StandsControl1_d_ct105_Image1" src="/stands.axd?image=DAVIVIENDA.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct106_h" href="/empresas-destacadas/trabajos-en-outsource_1259.aspx" >
                    <img id="StandsControl1_d_ct106_Image1" src="/stands.axd?image=logoStand-templateoutsource.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct107_h" href="/empresas-destacadas/trabajos-en-unicomer_1286.aspx" >
                    <img id="StandsControl1_d_ct107_Image1" src="/stands.axd?image=unicomer.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct108_h" href="/empresas-destacadas/trabajos-en-arqco_1595.aspx" >
                    <img id="StandsControl1_d_ct108_Image1" src="/stands.axd?image=t5f3bai1.vd4Arqco-principal.png" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct109_h" href="/empresas-destacadas/trabajos-en-banco-agricola_510.aspx" >
                    <img id="StandsControl1_d_ct109_Image1" src="/stands.axd?image=633632972816877070.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct110_h" href="/empresas-destacadas/trabajos-en-tigo_528.aspx" >
                    <img id="StandsControl1_d_ct110_Image1" src="/stands.axd?image=logo tigo.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct111_h" href="/empresas-destacadas/trabajos-en-banco-azteca_545.aspx" >
                    <img id="StandsControl1_d_ct111_Image1" src="/stands.axd?image=31l5gaoz.dv0Banco-azteca-principal.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct112_h" href="/empresas-destacadas/trabajos-en-consisa_558.aspx" >
                    <img id="StandsControl1_d_ct112_Image1" src="/stands.axd?image=50fyushd.hgaGrupo-consisa-principal-ajfsg.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct113_h" href="/empresas-destacadas/trabajos-en-banco-azul_1874.aspx" >
                    <img id="StandsControl1_d_ct113_Image1" src="/stands.axd?image=banco-azul-stand.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct114_h" href="/empresas-destacadas/trabajos-en-ria_1526.aspx" >
                    <img id="StandsControl1_d_ct114_Image1" src="/stands.axd?image=ria-stand1.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct115_h" href="/empresas-destacadas/trabajos-en-blanco-silva-consultoria-informatica_2171.aspx" >
                    <img id="StandsControl1_d_ct115_Image1" src="/stands.axd?image=wg3kdsvk.4fyBSCI-El-Salvador-principal.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct116_h" href="/empresas-destacadas/trabajos-en-omnisport_1254.aspx" >
                    <img id="StandsControl1_d_ct116_Image1" src="/stands.axd?image=logoStand-templateomnisport.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct117_h" href="/empresas-destacadas/trabajos-en-farmacias-economicas_1895.aspx" >
                    <img id="StandsControl1_d_ct117_Image1" src="/stands.axd?image=farmacias economicas logo.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct118_h" href="/empresas-destacadas/trabajos-en-mercosal_2395.aspx" >
                    <img id="StandsControl1_d_ct118_Image1" src="/stands.axd?image=njfhi4i1.3dplogo imagen mercosal.jpg" ></a>
            </span>
<span>
                <a id="StandsControl1_d_ct119_h" href="/empresas-destacadas/trabajos-en-hanes_570.aspx" >
                    <img id="StandsControl1_d_ct119_Image1" src="/stands.axd?image=hanesBoton.gif" ></a>
            </span>
    
    <span class="clear"></span>
</div>
<div id="nav-empresas">
    <a class="prev sprite-bkLink01" href="#">&lt;</a><a class="next sprite-bkLink01" href="#">&gt;</a>
</div>
    <a class="sprite-btnMedio sprite-btnMedio-align" href="/listado/empresas-destacadas.aspx">ver más empresas</a>
<span class="clear"></span>

                                    <span class="clear"></span>
                                </div>
                                <a id="s2_divTestimoniales" href="/empresas/testimoniales-de-empresas" target="_blank"><img id="s2_Image1" src="/Content/images/imgTestimonialesE.jpg" alt="Testimoniales de Empresas" style="border-width:0px;"></a>



    <div class="aliados">
        <div class="imgTitLanding-align sprite-imgTitLanding">
            nuestros aliados
        </div>
        <div class="contenido-landing">
            <p class="intro" style="text-align: justify;">
                Los siguientes medios anuncian nuestras ofertas de trabajo, comparten tips y te brindan informaci&oacute;n sobre nuestras iniciativas y ferias de trabajo ¡B&uacute;scalos!
            </p>
            <div class="panelesAliados">
                    <div class="aliado-item">
                        <a href="https://www.tecoloco.com.sv/MediaPartnersClick.ashx?mp=CvkgZs0bjgA%3d" class="partner-element" target="_blank">
                            <span class="partner">
                                <img class="partnerlogo" id="MediaPartnersControl1_DLMD_ctl00_Img" src="//content.tecoloco.com/Assets/mediapartner/aaeuhlb2.tdwLOGO_ZONAEMPLEO.jpg" style="width: 72px; height: 72px;">
                                Zona Empleo
                                <span class="clear"></span>
                            </span>
                        </a>
                    </div>
                    <div class="aliado-item">
                        <a href="https://www.tecoloco.com.sv/MediaPartnersClick.ashx?mp=mdy39hcMQs8%3d" class="partner-element" target="_blank">
                            <span class="partner">
                                <img class="partnerlogo" id="MediaPartnersControl1_DLMD_ctl00_Img" src="//content.tecoloco.com/Assets/mediapartner/rebw0lik.rtdLOGO_ELSALVADOR.COM.jpg" style="width: 72px; height: 72px;">
                                Elsalvador.com
                                <span class="clear"></span>
                            </span>
                        </a>
                    </div>
            </div>
            <div class="nav-aliados">
                <span class="nav-control"><a class="prev sprite-bkLink01" href="#">&lt;</a></span><span class="nav-control"><a class="next sprite-bkLink01" href="#">&gt;</a></span>
            </div>
            <span class="clear"></span>
        </div>
        <div class="foo-landing">
        </div>
    </div>
                            <span class="clear"></span>
                    </div>
                    


                        <meta name="keywords" content="trabajos en El Salvador, empleos en El Salvador, www.tecoloco.com.sv." />
    <meta name="description" content="Encuentra tu pr&#243;ximo trabajo hoy, las mejores ofertas de trabajo y ofertas de empleo en El Salvador con www.tecoloco.com.sv. Registrar tu curriculum en www.tecoloco.com.sv es gratis" />





<div class="hidden-desktop ">


    <div class="col-sm-12">

        <form action="/Default2.aspx" class="form-group">


            <div class="inner-addon left-addon">
                <i class="glyphicon glyphicon-search mobile-gris-oscuro"></i>



                <input class="Searchkeys form-control" id="Keywords" name="Keywords" onBlur="javascript:removeHtml(&#39;keysdektop&#39;);" onkeypress="javascript:stopRKey()" placeholder="Palabra clave" type="text" value="" />

            </div>
            <input class="btn btn-primary btn-only-tablet btnBuscarAhora" type="submit" name="s1$b1" id="s1_b1" value="Buscar ahora">
            <a class="btn btn-default btn-block btn-only-tablet" data-toggle="collapse" data-target="#filtrosBusqueda">Filtros de búsqueda</a>
            <span class="clear"></span>
            <div id="filtrosBusqueda" class="collapse">
                <select class="form-control categoria-dropdown" id="Categoria" name="Categoria"><option value="">Cualquier &#193;rea</option>
<option value="administrativo">Administraci&#243;n</option>
<option value="bodega-almacenamiento">Almacenamiento</option>
<option value="oficinas">Apoyo de Oficina</option>
<option value="banco-servicios-financieros">Banca | Servicios Financieros</option>
<option value="call-center">Call Center</option>
<option value="compras">Compras</option>
<option value="contabilidad">Finanzas | Contabilidad | Auditor&#237;a</option>
<option value="informatica-internet">Inform&#225;tica | Internet</option>
<option value="mantenimiento">Mantenimiento</option>
<option value="marketing-ventas">Mercadeo | Ventas</option>
<option value="logistica">Operaciones | Log&#237;stica</option>
<option value="ingenieria-calidad">Producci&#243;n | Ingenier&#237;a | Calidad</option>
<option value="publicidad">Publicidad | Comunicaciones | Servicios</option>
<option value="profesionales">Puestos Profesionales</option>
<option value="recursos-humanos">Recursos Humanos</option>
<option value="restaurantes">Restaurantes</option>
<option value="salud">Salud</option>
<option value="telefonia-telecomunicaciones">Telecomunicaciones</option>
<option value="otros-trabajos">Varios</option>
</select>
                <select class="form-control cargo-dropdown" id="Cargo" name="Cargo"><option value="">Cualquier Cargo</option>
</select>
                <select class="form-control" id="PaisId" name="PaisId"><option value="0">Centroam&#233;rica</option>
<option value="16">Costa Rica</option>
<option selected="selected" value="21">El Salvador</option>
<option value="29">Guatemala</option>
<option value="31">Honduras</option>
<option value="41">Nicaragua</option>
<option value="45">Panam&#225;</option>
<option value="53">Rep&#250;blica Dominicana</option>
</select>
                <input class="form-control" id="KeywordCompany" name="KeywordCompany" placeholder=" - compañía - " type="text" value="" />
                <span class="clear"></span>
            </div>
            <a class="btn btn-default btn-block btn-only-phone" data-toggle="collapse" data-target="#filtrosBusqueda">Filtros de búsqueda</a>
            <input class="btnBuscarAhora btn btn-primary btn-block btn-only-phone" type="submit" name="s1$b1" id="s1_b1" value="Buscar ahora">



            <span class="clear"></span>
        </form>


    </div>




    <span class="clear"></span>
</div>






<div class="mobile-content hidden-desktop">


    <h1 class="col-sm-12 col-xs-12">ofertas de trabajo, oportunidades de empleo </h1>


    
    <h2 class="col-sm-12 col-xs-12">&Uacute;ltimas ofertas publicadas</h2>

    <span class="clear"></span>

    <div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363449/vendedor-rutero.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=7550-636324236598876746.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Gestor de Cumplimiento (RUTA)</span>
            <br />
            
            Objetivo General: 
Validar el cumplimiento de preceptos relacionados con el man...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363449" data-job-title="Gestor de Cumplimiento (RUTA)" data-job-url="/363449/gestor-de-cumplimiento-ruta.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363449/vendedor-rutero.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363443/farmaceutico.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=635453571026562500.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >QU&#205;MICO DE LABORATORIO</span>
            <br />
            
            *Realizar análisis fisicoquímicso en las diferentes fases del proceso productivo...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363443" data-job-title="QU&#205;MICO DE LABORATORIO" data-job-url="/363443/quimico-de-laboratorio.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363443/farmaceutico.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-la-libertad"><i></i>La Libertad</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363437/disenador-grafico.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=40150-636548233406128562.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >OPERADOR DE PLOTTER</span>
            <br />
            
            OPERADOR DE PLOTTER DE IMPRESIÓN


DESCRIPCION DEL PUESTO:

Manejo de la má...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363437" data-job-title="OPERADOR DE PLOTTER" data-job-url="/363437/operador-de-plotter.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363437/disenador-grafico.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 23/03/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363433/chef.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=47980-636571351079655920.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Chef</span>
            <br />
            
            Realizar las preparaciones culinarias conforme a las recetas indicadas, empleand...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363433" data-job-title="Chef" data-job-url="/363433/chef.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363433/chef.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363432/medico.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=635458744369843750.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >MEDICO EMPRESARIAL</span>
            <br />
            
            Propósito:

Coordinar y dirigir el Sistema Médico de la planta por medio del e...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363432" data-job-title="MEDICO EMPRESARIAL" data-job-url="/363432/medico-empresarial.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363432/medico.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-la-libertad"><i></i>La Libertad</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363430/administrador.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=2633-636542245313808653.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Analista operativo</span>
            <br />
            
             Responsable administrativo del control  de solicitudes  enviadas a investigació...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363430" data-job-title="Analista operativo" data-job-url="/363430/analista-operativo.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363430/administrador.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363427/supervisor-de-mantenimiento.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=635127815946052500.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Coordinador  de Mantenimiento de Edificios e Insta...</span>
            <br />
            
            Empresa de Solido Prestigio desea contratar: Coordinador  de Mantenimiento de Ed...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363427" data-job-title="Coordinador  de Mantenimiento de Edificios e Instalaciones" data-job-url="/363427/coordinador-de-mantenimiento-de-edificios-e-instalaciones.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363427/supervisor-de-mantenimiento.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363408/asistente-contable.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=47916-636571359990724008.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Soporte de ventas Aviaci&#243;n</span>
            <br />
            
            Descripcion del puesto 
Administrar la facturación - precios de clientes de cré...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363408" data-job-title="Soporte de ventas Aviaci&#243;n " data-job-url="/363408/soporte-de-ventas-aviacion.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363408/asistente-contable.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 12/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363397/ejecutivo-de-ventas.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=635206408691588750.jpg" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >DEPENDIENTE DE SALA DE VENTAS SANTA TECLA Y ANTIGU...</span>
            <br />
            
            Grupo RAF

Requerimos contratar Señoritas
PLAZAS DISPONIBLES PARA: ANTIGUO CU...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363397" data-job-title="DEPENDIENTE DE SALA DE VENTAS SANTA TECLA Y ANTIGUO CUSCATLAN" data-job-url="/363397/dependiente-de-sala-de-ventas-santa-tecla-y-antiguo-cuscatlan.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363397/ejecutivo-de-ventas.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-la-libertad"><i></i>La Libertad</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div><div class="span12 plazaTablet tecoloco-wc">

    <div class="col-sm-10 col-xs-10 mobile-plaza-content">



        <a href="/363364/ejecutivo-pyme.aspx?fromApp=true" class="mobile-job-link" >
            
            <img src="/logo.axd?image=2618-635811980646571320.png" alt="" style="height: 100px; width: 100px;" class="logo thumbnail" />            
            
            <span class="mobile-job-name" >Ejecutivo PYME</span>
            <br />
            
            Ejecutivo PYME
San Salvador

Objetivo de Puesto:
Promover los productos dest...
            <span class="clear" ></span>
        </a>
       
    </div>
    <div class="col-sm-2 col-xs-2 btn-container dropdown">
        <a class="btn-menu dropdown-toggle" data-toggle="dropdown"></a>
        <ul class="dropdown-menu dropdown-menu-right">

            

                <li>



                        <a style="cursor: pointer;" class="save-job job-btn floatR btnAplica" data-jobid="363364" data-job-title="Ejecutivo PYME" data-job-url="/363364/ejecutivo-pyme.aspx">
                            <span class="saved mleft5 mtop3"></span><span class="data-location-txt"><i></i>Agregar como favorito</span>
                        </a>

                </li>
            <li class="divider"></li>

            
                <li>
                    <a class="verOferta" href="/363364/ejecutivo-pyme.aspx"  style="cursor: auto;"><i></i>Ver oferta</a>
                </li>

            <li class="divider"></li>
            
            <li>
                <span>Fecha fin: 19/04/2018</span>
            </li>


                <li><span>El Salvador</span></li>
                        <li><a href="/trabajos-en-san-salvador"><i></i>San Salvador</a></li>

        </ul>
    </div>



    <span class="clear"></span>






</div>

    <span class="clear"></span>
</div>



<div class="mainContent visible-desktop">

    
    <form action="/Default2.aspx" method="GET">
        
        <div class="sprite-bkBusqueda-align sprite-bkBusqueda barG">
            <h2>caja de búsqueda de trabajo</h2>
            <span class="clear"></span>
            <span class="inputText areas">
                <select class="span12 categoria-dropdown" id="Categoria" name="Categoria"><option value="">Cualquier &#193;rea</option>
<option value="administrativo">Administraci&#243;n</option>
<option value="bodega-almacenamiento">Almacenamiento</option>
<option value="oficinas">Apoyo de Oficina</option>
<option value="banco-servicios-financieros">Banca | Servicios Financieros</option>
<option value="call-center">Call Center</option>
<option value="compras">Compras</option>
<option value="contabilidad">Finanzas | Contabilidad | Auditor&#237;a</option>
<option value="informatica-internet">Inform&#225;tica | Internet</option>
<option value="mantenimiento">Mantenimiento</option>
<option value="marketing-ventas">Mercadeo | Ventas</option>
<option value="logistica">Operaciones | Log&#237;stica</option>
<option value="ingenieria-calidad">Producci&#243;n | Ingenier&#237;a | Calidad</option>
<option value="publicidad">Publicidad | Comunicaciones | Servicios</option>
<option value="profesionales">Puestos Profesionales</option>
<option value="recursos-humanos">Recursos Humanos</option>
<option value="restaurantes">Restaurantes</option>
<option value="salud">Salud</option>
<option value="telefonia-telecomunicaciones">Telecomunicaciones</option>
<option value="otros-trabajos">Varios</option>
</select>


            </span>
            <span class="inputText cargos">
                <select class="span12 cargo-dropdown" id="Cargo" name="Cargo"><option value="">Cualquier Cargo</option>
</select>
                
            </span>
            <span class="inputText paises">
                <select class="span12" id="PaisId" name="PaisId"><option value="0">Centroam&#233;rica</option>
<option value="16">Costa Rica</option>
<option selected="selected" value="21">El Salvador</option>
<option value="29">Guatemala</option>
<option value="31">Honduras</option>
<option value="41">Nicaragua</option>
<option value="45">Panam&#225;</option>
<option value="53">Rep&#250;blica Dominicana</option>
</select>
                
            </span>

            <span class="inputText compania">
                <input id="KeywordCompany" name="KeywordCompany" placeholder="introduce el nombre de una compañía" type="text" value="" />
            </span>

            <span class="inputText busqueda">
                <input class="Searchkeys keysmovil" id="Keywords" name="Keywords" onBlur="javascript:removeHtml(&#39;keysmovil&#39;);" onkeypress="javascript:stopRKey()" type="text" value="" />
                
                <button class="btnBusquedaBox-align sprite-btnBusquedaBox" name="s1$b1" id="s1_b1" value=""></button>
            </span>
        </div>
    </form>

    <div>
        

        <div class="sprite-bkListadoOfertas-align sprite-bkListadoOfertas visible-desktop">
            <h1>ofertas de trabajo, oportunidades de empleo</h1>
            <h2>últimas ofertas publicadas</h2>
        </div>
        <div style="padding: 0 22px;">
            <span class="plaza visible-desktop">
    <img  src="/logo.axd?image=7550-636324236598876746.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363449/vendedor-rutero.aspx"  style="cursor: auto;">Gestor de Cumplimiento (RUTA)</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        Objetivo General: 
Validar el cumplimiento de preceptos relacionados con el manejo de inventarios, cartera y efectivo por los encargados de ruteo del área comercial, con base a los controles acordados con la D... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363449/vendedor-rutero.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363449" data-job-title="Gestor de Cumplimiento (RUTA)" data-job-url="/363449/gestor-de-cumplimiento-ruta.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=635453571026562500.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363443/farmaceutico.aspx"  style="cursor: auto;">QU&#205;MICO DE LABORATORIO</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-la-libertad" class="lugar-trabajo">La Libertad</a>
    
    <span class="detalle-trabajo">
        *Realizar análisis fisicoquímicso en las diferentes fases del proceso productivo, procurando se lleven a cabo en los tiempos definidos y garantizando la confiabilidad de los resultados, de acuerdo con normas y ... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363443/farmaceutico.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363443" data-job-title="QU&#205;MICO DE LABORATORIO" data-job-url="/363443/quimico-de-laboratorio.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=40150-636548233406128562.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363437/disenador-grafico.aspx"  style="cursor: auto;">OPERADOR DE PLOTTER</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        OPERADOR DE PLOTTER DE IMPRESIÓN


DESCRIPCION DEL PUESTO:

Manejo de la máquina de impresión y encargado de las muestras de color.

REQUISITOS: 

•	Edad: mínima 22 años a 40 años
•	Nivel Académico: G... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />23/03/2018</span>
        <a class="verOferta" href="/363437/disenador-grafico.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363437" data-job-title="OPERADOR DE PLOTTER" data-job-url="/363437/operador-de-plotter.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=47980-636571351079655920.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363433/chef.aspx"  style="cursor: auto;">Chef</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        Realizar las preparaciones culinarias conforme a las recetas indicadas, empleando las técnicas, tipo, calidad y cantidad de ingredientes requeridos, así como los equipos y utensilios, con base en los estándares... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363433/chef.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363433" data-job-title="Chef" data-job-url="/363433/chef.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=635458744369843750.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363432/medico.aspx"  style="cursor: auto;">MEDICO EMPRESARIAL</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-la-libertad" class="lugar-trabajo">La Libertad</a>
    
    <span class="detalle-trabajo">
        Propósito:

Coordinar y dirigir el Sistema Médico de la planta por medio del establecimiento de Políticas y Procedimientos de un sistema de servicio médico completo y que a la vez gestione medidas de salud pr... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363432/medico.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363432" data-job-title="MEDICO EMPRESARIAL" data-job-url="/363432/medico-empresarial.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=2633-636542245313808653.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363430/administrador.aspx"  style="cursor: auto;">Analista operativo</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
         Responsable administrativo del control  de solicitudes  enviadas a investigación por los Jefes Validadores de Crédito, generación de reportes relacionados con los diferentes estatus de dichas solicitudes, segu... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363430/administrador.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363430" data-job-title="Analista operativo" data-job-url="/363430/analista-operativo.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=635127815946052500.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363427/supervisor-de-mantenimiento.aspx"  style="cursor: auto;">Coordinador  de Mantenimiento de Edificios e Instalaciones</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        Empresa de Solido Prestigio desea contratar: Coordinador  de Mantenimiento de Edificios e Instalaciones

Requisitos:
*Edad: 25 a 45 años.
*Nivel académico: Egresado de Arquitectura.(Indispensable)
*Experie... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363427/supervisor-de-mantenimiento.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363427" data-job-title="Coordinador  de Mantenimiento de Edificios e Instalaciones" data-job-url="/363427/coordinador-de-mantenimiento-de-edificios-e-instalaciones.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=47916-636571359990724008.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363408/asistente-contable.aspx"  style="cursor: auto;">Soporte de ventas Aviaci&#243;n </a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        Descripcion del puesto 
Administrar la facturación - precios de clientes de crédito.

Requisitos:
1. Bilingue
2. Experiencia de 2 años como auxiliar administrativo - contable
3. Manejo de paquete de Ofimá... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />12/04/2018</span>
        <a class="verOferta" href="/363408/asistente-contable.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363408" data-job-title="Soporte de ventas Aviaci&#243;n " data-job-url="/363408/soporte-de-ventas-aviacion.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=635206408691588750.jpg" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363397/ejecutivo-de-ventas.aspx"  style="cursor: auto;">DEPENDIENTE DE SALA DE VENTAS SANTA TECLA Y ANTIGUO CUSCATLAN</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-la-libertad" class="lugar-trabajo">La Libertad</a>
    
    <span class="detalle-trabajo">
        Grupo RAF

Requerimos contratar Señoritas
PLAZAS DISPONIBLES PARA: ANTIGUO CUSCATLAN Y SANTA TECLA

COMPETENCIAS REQUERIDAS:
- Conocimientos de tecnológicos, computación y ventas
-Pro activa 
-Excelente... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363397/ejecutivo-de-ventas.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363397" data-job-title="DEPENDIENTE DE SALA DE VENTAS SANTA TECLA Y ANTIGUO CUSCATLAN" data-job-url="/363397/dependiente-de-sala-de-ventas-santa-tecla-y-antiguo-cuscatlan.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>




<span class="plaza visible-desktop">
    <img  src="/logo.axd?image=2618-635811980646571320.png" alt="" style="height: 100px; width: 100px;" class="logo" />
            
           <a class="oferta-trabajo" href="/363364/ejecutivo-pyme.aspx"  style="cursor: auto;">Ejecutivo PYME</a>
    
    
   
            <span class="pais-trabajo" >El Salvador</span>
                <a href="/trabajos-en-san-salvador" class="lugar-trabajo">San Salvador</a>
    
    <span class="detalle-trabajo">
        Ejecutivo PYME
San Salvador

Objetivo de Puesto:
Promover los productos destinados a la Pequeña y Mediana Empresa. Administrar la cartera de clientes con este perfil con base en la estrategia de negocios y ... 
    </span>    
    <span class="imgVigencia-align sprite-imgVigencia">
        Fecha fin<br />19/04/2018</span>
        <a class="verOferta" href="/363364/ejecutivo-pyme.aspx" target="_blank" style="cursor: auto;">Ver oferta</a>
    
            <a class="save-job agregar-oferta-favorito " data-jobid="363364" data-job-title="Ejecutivo PYME" data-job-url="/363364/ejecutivo-pyme.aspx" onclick="var s=s_gi(&#39;stepstone-saongroup-tecoloco-prod&#39;);s.linkTrackVars=&#39;events,props,server,evars&#39;;s.linkTrackEvents =&#39;event16&#39; ;s.events=&#39;event16&#39; ;s.tl(this,&#39;o&#39;,&#39;listing save&#39;);" >
                <span class="saved"></span><span class="data-location-txt">Agregar como favorito</span>
            </a>
    
    <span class="clear"></span>
</span>
<br />
<span class="clear"></span>





        </div>


        


        

        <!-- TecoAds_468_15_2013_2 -->
        

    </div>
</div>

<script type="text/javascript">
    var stopSubmit = false;

    function stopRKey(evt) {
        evt = (evt) ? evt : ((event) ? event : null);
        var node = (evt.target) ? evt.target : ((evt.srcElement) ? evt.srcElement : null);
        if ((evt.keyCode == 13) && (node.type == "text")) {
            stopSubmit = true;
            return false;
        }
        stopSubmit = false;
        return true;
    }

    $(function () {


        $(".Searchkeys").keyup(function() {
            var str = $(this).val();
            if (/[~`!#$%\^&*+=\-\[\]\\';,/{}|\\":<>\?]/g.test(str)) {
                $('.btnBuscarAhora').attr("disabled", "disabled");
                $(".Searchkeys").addClass("ErrorTextBox");
                $(".btnBuscarAhora").attr("title", "Ha ingresado caracteres no permitidos");

                //alert('Caracteres no permitidos');

                //str = str.replace(/<[\/]{0,1}([A-Z]|[a-z])[^><]*>/g, '');
                //str = str.replace(/&nbsp;/g, '');
                //str = str.replace(/'/g, '');
                //var txt = str;
                //$('.btnBuscarAhora').val(txt);
                stopSubmit = true;
                return false;
            } else {
                $(".Searchkeys").removeClass("ErrorTextBox");
                $(".btnBuscarAhora").attr("title", "Buscar");
                $('.btnBuscarAhora').removeAttr("disabled");
                stopSubmit = false;
                return true;
            }
        });

        $(".categoria-dropdown").change(function() {
            $.ajax({ url: "/Jobs/GetCargos", data: { area: $(this).find("option:selected").text() } }).success(function(data) {
                $('.cargo-dropdown').html('');
                $.each(data, function(i, value) {

                    $('.cargo-dropdown').append($('<option>').text(value.Description).attr('value', value.Id));
                });
            });

        });

        $("form").submit(function(e) {
            if (stopSubmit) {
                e.preventDefault();
                stopSubmit = false;
                return false;
            } else {
                return true;
            }
        });

    });

    function removeHtml(id) {
        var str = $("." + id).val();
        if (/[~`!#$%\^&*+=\-\[\]\\';,/{}|\\":<>\?]/g.test(str)) {
            alert('Caracteres no permitidos');
            str = str.replace(/<[\/]{0,1}([A-Z]|[a-z])[^><]*>/g, '');
            str = str.replace(/&nbsp;/g, '');
            str = str.replace(/'/g, '');
            var txt = str;
            $("." + id).val(txt);
            return false;
        } else {
            return true;
        }
    };

</script>

<div id="modal_newcv" class="modal fade" role="dialog">
    <div class="modal-dialog">
        <!-- Modal content-->
        <div class="modal-content">
            <div class="modal-header">
                <a class="close" data-dismiss="modal">&times;</a>
                <h4 class="modal-title">NUEVO CURRÍCULO</h4>
            </div>
            <div class="modal-body">
                <div id="wrap_Experiencias">
                    
<div id="NewCurriculum" title="Crear Nuevo Curriculum" class="tecoModal">
    <div class="panel-oferta trabajo-formulario edicion" style="border: none;">
        <div class="left-TA visible-sm-inline col-sm-2">
            <span class="txRed">*</span>
            <span class="visible-lg-inline">T&iacute;tulo o nombre de curr&iacute;culum:</span>
            <span class="visible-sm-inline hidden-desktop">T&iacute;tulo de curr&iacute;culum:</span>
        </div>
        <div class="right-TA col-sm-10 col-xs-12">
            <input type="text" maxlength="50" id="txt_titlecv" class="form-control" placeholder="T&iacute;tulo o nombre de curr&iacute;culum">
            <br class="visible-desktop">
            <span style="color:Red;display:none; font-size: 11px;">(*) requerido</span>
            <br class="visible-desktop">
            <div id="ctl00_CP_rlstTipo">
                <input type="radio" name="CvTipo" value="1" checked="checked"> P&uacute;blico
                <input type="radio" name="CvTipo" value="0"> Privado
            </div>
        </div>
        <br class="visible-desktop">
        <br class="visible-desktop">

        <div class="linePun visible-desktop">
        </div>


        <span class="clear"></span>
        <span class="sep visible-desktop"></span>
        <br />

        <a class="hidden-desktop btn btn-default btn-block btnDrop" data-toggle="collapse" data-target="#panel_des">Descripciones de tipos<span class="caret"></span></a>


        <p id="panel_des" class="col-md-12 col-xs-12m m-t-10 collapse">


            <span class="txRed red">
                Público:
            </span>
            <br>
            <span class="txt-informativo-normal">
                Cuando tu curr&iacute;culum sea consultado por una empresa esta podrá visualizar todos los datos del mismo.
            </span>
            <br>
            <span class="txRed red">
                Privado:
            </span>
            <br>
            <span class="clear"></span>
            <span class="txt-informativo-normal">
                Cuando tu curr&iacute;culum sea consultado por una empresa no se podrá visualizar tu nombre y tu actual lugar de trabajo.
            </span>
            <span class="clear"></span>

            <br class="visible-desktop" /><br />
        </p>
        
        
        
        <br/>

        <a id="ctl00_CP_defaultBtn" class="btnAplica floatL btn btn-primary col-xs-5 col-sm-5 visible-phone" href="#" onclick="javascript:saveCV();" style="margin-top: 5px;">Guardar</a>
        <a class="btnAplica floatL btn btn-primary col-xs-5 col-xs-offset-2 col-sm-offset-2 col-sm-5 visible-phone" href="#" onclick="javascript:closeNewCv();" data-dismiss="modal" style="margin-top: 5px;">Cancelar</a>

        <a id="ctl00_CP_defaultBtn" class="btnAplica floatL visible-desktop" href="#" onclick="javascript:saveCV();" style="margin-top: 5px;">Guardar</a>
        <a class="btnAplica floatL visible-desktop" href="#" onclick="javascript:closeNewCv();" data-dismiss="modal" style="margin-top: 5px;">Cancelar</a>

        <span class="clear"></span>
    </div>

</div>
                </div>
            </div>
            <div class="modal-footer">
                
            </div>
        </div>

    </div>
</div>


<script src="/Scripts/aliados.js" type="text/javascript"></script>





                    

                    <span class="clearfix"></span>

                </div>
            </div>






<link href="/Content/estilosprite.css" media='screen and (min-width: 1024px)' rel="stylesheet" />

<div class="foo hidden-phone">
    <div class="content row-fluid">
        <div class="span12 left">
            <div class="pl">
                <p>Descarga nuestra app, disponible en:</p>







                <ul>

                    <li class="pull-left"><a href="https://itunes.apple.com/us/app/tecoloco.com-bolsa-trabajo/id1134960846" target="_blank"><img src="/Content/images/appStore.png" alt="App Store" /></a></li>
                    <li class="pull-left"><a href="https://play.google.com/store/apps/details?id=com.stepstone.tecoloco&amp;hl=es" target="_blank"><img src="/Content/images/googlePlay.png" alt="Google Play" /></a></li>

                </ul>
                    
                <span class="clear"></span>


                    <span class="titFoo">© Tecoloco.com</span>    
                <br />

                <span class="anyo">2013 </span>Todos los Derechos Reservados<br>
                <span class="visible-desktop">
                    Esta página esta optimizada para: <a href="https://www.mozilla-europe.org/es/firefox/" rel="nofollow" target="_blank" class="txLine txB">Firefox 3.5+ </a>,<a href="https://www.microsoft.com/es-es/download/internet-explorer.aspx" rel="nofollow" target="_blank" class="txLine txB"> Internet Explorer 8+ </a>,<a href="https://www.google.com/chrome/" rel="nofollow" target="_blank" class="txLine txB"> Google Chrome </a>
                    <br>
                </span>
                <br>
                |<a href="/ ">Inicio</a>
                |
 <a id="SM_l4" href="/default2.aspx">Búsqueda de Empleos</a>                 |
                
 <a href="/contacto.aspx">Contáctanos</a>                 |
                
 <a href="/frmFeed.aspx">Rss Feed</a>                 |

                
 <a href="/frmQSomos.aspx">Quienes Somos</a>                 |

                <span class="visible-desktop">

                
                
                
                
                    

 <a href="/frmPreguntas.aspx">Preguntas</a>                |
                <a id="SM_l11" href="/Empresas/registro_empresa1.aspx">Registro Empresas</a>
                |
  <a id="SM_l12" href="/Candidatos/frmAbreCuenta.aspx">Registro Candidatos</a>                    
                |
 <a id="SM_l13" href="/SiteMaps.aspx">Mapa del Sitio</a>                 <br />
                |
                
                <a href="/login.aspx">Ingreso Candidatos</a>
                |

                <a id="SM_l15" href="/loginEmpresas.aspx">Ingreso Empresas</a>


                <span id="SM_SpanSugerencias">
                    |<a id="SM_l16" href="mailto:info@tecoloco.com">Sugerencias</a>
                </span>
                
                |
                
                    
                    <a href="/empresas.aspx">Directorios de Empresas</a>  
                |
                    


                    
                        <a id="SM_HyperLink1" href="/tecoAds/frmCreateAds.aspx">Anuncios con Tecoloco</a> |
                    
                
                    
                        <a id="SM_hlblog" href="/Blog" target="_self">Blog</a> |    
                <a href="/thenetwork.aspx">Reclutamiento Internacional</a>
                </span>
            </div>
            <div class="pr hidden-phone">

                <div class="redes">
 <a id="SM_ShortCuts1_rsslink" class="sprite-btnRss" rel="nofollow" href="/frmfeed.aspx" target="_self"></a>                    <a id="SM_ShortCuts1_lnkYouTube" class="sprite-btnYouTube" rel="nofollow" href="https://www.youtube.com/user/TecolocoSupport/" target="_blank"></a>
                    <a id="SM_ShortCuts1_lnkTwitter" class="sprite-btnTwitter" rel="nofollow" href="https://twitter.com/TrabajosSV" target="_blank"></a>
                    <a id="SM_ShortCuts1_lnkFacebook" class="sprite-btnFB" rel="nofollow" href="https://www.facebook.com/EmpleoElSalvador" target="_blank"></a>
                    <a id="SM_ShortCuts1_lnkG" class="sprite-btnG" rel="nofollow" href="https://plus.google.com/+TecolocoSv" target="_blank"></a>
                    <a id="SM_ShortCuts1_lnkLkdIn" class="sprite-btnLinkedInRS" rel="nofollow" href="https://www.linkedin.com/company/tecoloco-com" target="_blank"></a>

                        <a id="SM_ShortCuts1_HyperLink2" class="sprite-btnBlogRS" href="https://www.tecoloco.com.sv/blog" target="_self"></a>

                    

                </div>
 <img id="SM_fooLogo" class="logoFoo" src="/Content/images/logoTecolocoFoo.jpg" style="border-width: 0px;">                <div class="saon">
                    <span class="titFoo">Una empresa de:</span>
                    <br>
                    <a id="SM_Image2" class="logoFoo sprite-logoSaonGroup" style="border-width: 0px;" href="https://saongroup.com/" target="_blank">
                        
                        </a>
                </div>
            </div>
        </div>
    </div>
</div>

<div class="phone visible-phone foo appstore">

    <p class="col-xs-12 col-sm-12">Descarga nuestra app, disponible en:</p>

    <ul class="list-unstyled">

        <li class="pull-left"><a href="https://itunes.apple.com/us/app/tecoloco.com-bolsa-trabajo/id1134960846" target="_blank"><img src="/Content/images/appStore.png" alt="App Store" /></a></li>
        <li class="pull-left"><a href="https://play.google.com/store/apps/details?id=com.stepstone.tecoloco&amp;hl=es" target="_blank"><img src="/Content/images/googlePlay.png" alt="Google Play" /></a></li>

    </ul>

    <span class="clear"></span>

 <span>© Tecoloco.com</span>     <span class="anyo">2013 </span>Todos los Derechos Reservados<br><br>

    <span class="clear" ></span>

                <a href="/" >Inicio</a>
                
 <a href="/default2.aspx">Búsqueda de Empleos</a>                 

 <a href="/contacto.aspx">Contáctanos</a>      

 <a href="/frmFeed.aspx">Rss Feed</a>                 


 <a href="/frmQSomos.aspx">Quienes Somos</a>                 


    
    
    
    
 <a href="/frmPreguntas.aspx">Preguntas</a>    
    
    
  <a href="/Candidatos/frmAbreCuenta.aspx">Registro Candidatos</a> 
    
 <a href="/SiteMaps.aspx">Mapa del Sitio</a>     
    
    <a href="/login.aspx">Ingreso Candidatos</a>
    

    

    
    
        <a href="mailto:info@tecoloco.com">Sugerencias</a>
    

    <a href="/empresas.aspx">Directorios de Empresas</a>
    


    

    
        <a id="SM_hlblog" href="/Blog" target="_self">Blog</a>


        
    <div class="productVersion" style="width: 90%; height: 40px; background-color: white; margin:auto; padding: 10px; display: none;">
        Environment: www.tecoloco.com.sv, Build Version: V 1.0.0.0, Date Release: 09/03/2018
    </div>

    <span class="clear" ></span>

</div>

            <div id="session">
                <ul>
                    <li class="user">
                        <a title="Ingresa a tu cuenta" class="tt" href="/login.aspx">
                                <img id="ctl00_LoginCandidato1_imgFoto" src="/Content/images/nopicuser.jpg" />
                        </a>
                        <a title="Ingresa a tu cuenta" class="tt" href="/login.aspx">
                            <span>Mi Cuenta:</span>
                        </a>
                        <br />
                        <!--:::::: USERNAME ::::::
                    si no existe nada dentro de este link (que tiene la clase username) entonces
                    aparecerán los links para registrarse e iniciar sesión automáticamente-->



                        <a title="Ingresa a tu cuenta" class="username tt" href="/Candidate"></a>



                        <!--:::::: FIN USERNAME ::::::-->
                        <br />
                        <a class="cerrar" href="/logout">-cerrar sesión-</a>
                    </li>
                    <!--::::::::::::::::: CURRICULOS :::::::::::::::::::::::::::
                Esta es la estructura de los currículo almacenados del candidato
                cada div con la clase "cv" es una estructura de currículo-->

                    <li class="cvs">
                        <div class="misCvs">
                            <div class="wrapCvs visible-desktop">
                                <!--::::::::::::::::: FIN CURRICULOS :::::::::::::::::::::::::::-->
                                <!--                    ::::::::::::::::::: BOTON DE REGISTRO DE CV'S :::::::::::::::::::::::
                            Si no esxiste ni un div con la clase "cv" este botón aparecerá para que el candidato
                            vaya directamente a registrar su o sus currículos-->
                                <div class="registraCV">
                                    <a href="javascript:addNewCv();" class="sprite-btnRegistroCvUser">
                                        
                                    </a>
                                </div>
                                <!--                    ::::::::::::::::::: BOTON DE REGISTRO DE CV'S :::::::::::::::::::::::  -->

                            </div>
                        </div>
                        <div class="visible-desktop">
                            <div class="barra ">
                            </div>
                            <span class="completado">completado</span>
                            <a href="#" class="nextCV sprite-btnNextCv">
                                
                            </a>
                            <a href="#" class="prevCV sprite-btnPrevCv">
                                
                            </a>
                        </div>
                    </li>
                </ul>
                <div class="visible-desktop">
                    <div class="medidor">
                        <span class="numero"></span>
                    </div>
                    <a href="#" class="userHelp verAyuda sprite-btnUserHelp" title="AYUDA del panel de CV's:&lt;br/&gt;&lt;br /&gt;Muestra información relevante de tu(s) currículo(s) almacenado(s) en tu cuenta.&lt;br /&gt;&lt;br /&gt;ACCIONES:&lt;br/&gt;&lt;br/&gt;BOTÓN ACTUALIZAR: Utilízalo para refrescar la fecha de actualización de tu CV (sin modificar información).&lt;br /&gt;&lt;br /&gt;BOTÓN EDITAR: Utilízalo para modificar la información de tu CV." style="display: block;">
                        
                    </a>
                </div>
            </div>
            <div id="contenedor-ayuda">
                <div class="logoAyuda">
                </div>
                <span class="contenido-ayuda"></span>
            </div>
            <div id="contenedor-tooltip">
            </div>
            <div style="display: none;">
               
            </div>
            <script type="text/javascript">
    $(function () {
        //$("#NewCurriculum").dialog({ autoOpen: false, width: 600, modal: true });
        //$('#modal_newcv').modal('show');
    });

    $(document).ready(function () {
        $(".save-job").live('click', function () {
                        
            var cookieName = 'saved_jobs';
            var jobId = $(this).data('jobid');
            var jobTitle = $(this).data('job-title');
            var jobIds;
            
            if (!$.cookie(cookieName)) {
                $.cookie(cookieName, JSON.stringify([{ id: jobId, title: jobTitle }]), { path: '/' });
            } else {
                jobIds = JSON.parse($.cookie(cookieName), { path: '/' });
                jobIds.unshift({ id: jobId, title: jobTitle });
                $.cookie(cookieName, JSON.stringify(jobIds), { path: '/' });
            }
            $(this).addClass('save-job agregar-oferta-favorito job-saved');
            $(this).children(".data-location-txt").html("Agregado a favoritos");
            showNotification("La oferta se guardará en tus Ofertas Almacenadas la próxima vez que inicies sesión.<a href=\"/login.aspx\"> Ir a inicio de sesión</a>");
            


        });

    });

    function addNewCv() {
        //$('#NewCurriculum').dialog('open');
        $('#modal_newcv').modal('show');
    }

    function closeNewCv() {
        //$('#NewCurriculum').dialog('close');
        $('#modal_newcv').modal('hide');
    }

    function saveCV() {
        if (window.grecaptcha.getResponse().length === 0) {
            $("#recaptcha-error-div").addClass("recaptcha-error");
            $("#recaptcha-error-message-div").html("Comprueba que no eres un robot.");
            return;
        }

        if ($("input[name='CvTipo']:checked").val() != "undefined" && $("#txt_titlecv").val() != "") {
            $.ajax({
                url: "/Curriculum/SaveNameAndType",
                type: 'POST',
                data: ko.toJSON({ 
                    id: "0",
                    name: $("#txt_titlecv").val(), 
                    isPublic: ($("input[name='CvTipo']:checked").val()=="1")
                    ,recaptchaCode: grecaptcha.getResponse()
                }),
                dataType: "json",
                contentType: 'application/json; charset=utf-8',
                success: function(newCvId) {
                    if (newCvId != null) {
                        window.location.href = '/Candidato/Curriculum/Edit?id=' + newCvId;
                        //$("#NewCurriculum").dialog("close");
                    }
                    else {
                        alert("Ocurrió un problema almacenando los datos, por favor intente nuevamente");
                        grecaptcha.reset();
                    }
                }
            });
        } else {
            alert("Debe completar los campos");
        }

    }
            </script>

            
<div id="btn_feedback">
    
    <a href="javascript:getFeedData();" class="sprite-feedback-align sprite-feedback"></a>
</div>




<div id="modal_feedback" class="modal fade" role="dialog">
    <div class="modal-dialog">

        <!-- Modal content-->
        <div class="modal-content">
            <div class="modal-header">
                <button type="button" class="close" data-dismiss="modal">&times;</button>
                <h4 class="modal-title">Sugerencias</h4>
            </div>
            <div class="modal-body">
                
                
                
                
                <div id="div_feedback" class="floatL recentsearch-txt hide">

                    <div class="left-TA" >
                        <label class="left">Nombre: </label>
                    </div>
                    <div class="right-TA" >
                        <input class="form-control feed_controls" type="text" id="txt_namefeed" style="" />
                    </div>
                    <div class="clear"></div>
                    <br />
                    <div class="left-TA">
                        <label class="Profile_Title">(*)Email: </label>
                    </div>
                    <div class="right-TA">
                        <input class="form-control feed_controls" type="text" id="txt_emailfeed" /><label id="lb_valmailfeed" class="required-field">Campo Requerido</label>
                    </div>
                    <div class="clear"></div>
                    <br />
                    <div class="right-TA" >
                        <label class="Profile_Title">(*)Mensaje:</label>
                    </div>
                    
                    
                    <textarea maxlength="2000" id="txt_messagefeed" class="form-control feed_controls" ></textarea>
                    
                    <label id="lb_valmessagefeed" class="required-field">Campo requerido</label>
                    <div class="clear"></div>
                    <br />
                    <span class="clear"></span>
                    <div class="floatR">
                        
                    </div>


                </div>



            </div>
            <div class="modal-footer">
                <button type="button" class="btn btn-default"  onclick="javascript:PostFeedback(); ">Enviar</button>
                <button type="button" class="btn btn-default"  onclick="javascript:CloseFeedBack(); ">Cerrar</button>
            </div>
        </div>

    </div>
</div>







<script type="text/javascript">
    
    function getFeedData() {
        $.ajax({
            cache: false,
            url: "/Home/GetDataFeedBack",
            type: 'Get',
            contentType: 'application/json; charset=utf-8',
            success: function (data) {
                if (data != null) {
                    $("#txt_namefeed").val(data.name);
                    $("#txt_emailfeed").val(data.mail);




                    //$("#div_feedback").data("kendoWindow").open().center();
                    $('#modal_feedback').modal('show');







                } else {
                    $("#txt_namefeed").val("");
                    $("#txt_messagefeed").val("");
                    $("#txt_emailfeed").val("");
                }
            }
        });
    }

    $(function () {
        $("#div_feedback").removeClass("hide");
        $("#lb_valmailfeed").hide();
        $("#lb_valmessagefeed").hide();
        




        //$("#div_feedback").kendoWindow({ width: '550px', title: 'SUGERENCIAS', modal: true, visible: false, position: ['center', 'center'] });
        //$('#modal_feedback').modal('show');



    });

    function PostFeedback() {
        var url = "";
        if ($("#txt_emailfeed").val() == "")
            $("#lb_valmailfeed").show();
        if ($("#txt_messagefeed").val() == "")
            $("#lb_valmessagefeed").show();
        if ($("#txt_emailfeed").val() != "" && $("#txt_messagefeed").val() != "") {
            $.ajax({
                url: '/Home/PostFeedback',
                type: 'POST',
                data: { name: $("#txt_namefeed").val(), message: $("#txt_messagefeed").val(), email: $("#txt_emailfeed").val(), url: url },
                success: function (data) {
                    if (data == "1") {
                        alert("Sugerencia enviada satisfactoriamente.");






                        //$("#div_feedback").data("kendoWindow").close();
                        $('#modal_feedback').modal('hide');





                        $("#txt_namefeed").val("");
                        $("#txt_messagefeed").val("");
                        $("#txt_emailfeed").val("");
                        $("#lb_valmailfeed").hide();
                        $("#lb_valmessagefeed").hide();
                    } else if (data == "2") {
                        alert("Sugerencia no enviada, favor intentar nuevamente.");
                    } else {
                        alert("Error al enviar tu sugerencia, " + data);
                    }
                }
            });
        }

    }

    function CloseFeedBack() {
        $("#txt_namefeed").val("");
        $("#txt_messagefeed").val("");
        $("#txt_emailfeed").val("");
        $("#lb_valmailfeed").hide();
        $("#lb_valmessagefeed").hide();





        //$("#div_feedback").data("kendoWindow").close();
        $('#modal_feedback').modal('hide');
    }
</script>

            
            

            

            <div id="sticky-notification" style="display: none;" class="fixedNotif z-notif">
                <div id="notif">
                    <div id="full-notif">
                        


    <div id="notification" class="DashboardNotificationBox" style="float: left; position:relative;">
        <div>






            <div id="notificationIcon"></div>
            
            <div class="dashgray-txt message"s></div>            
            
            <div id="closeNotification"><div id="closeNotificationIcon"></div></div> 




        </div>
        </div>

                    </div>
                </div>
            </div>
                <script type="text/javascript">
        var report_suite_id = 'stepstone-saongroup-tecoloco-prod';
    </script>
    <script src="/Scripts/VisitorAPI.js"></script>
    <script src="/Scripts/AppMeasurement.js"></script>
    <script language="JavaScript" type="text/javascript">
        s.account = report_suite_id;



        s.prop1 = "";
        s.prop4 = "";
        s.prop6 = "SV";
        s.prop7 = "ES";
        s.prop9 = "";
        s.prop10 = "";
        s.prop11 = "";
        s.prop28 = "CCBot/2.0 (http://commoncrawl.org/faq/)";
        s.prop35 ="https://www.tecoloco.com.sv/";
        s.prop36 = "1.2.1";
        s.channel = "Home Page";
        s.pageName = "Home Page";
        s.server = "www.tecoloco.com.sv";
        s.eVar15 = s.server;
        s.hier1 = s.prop6 + ":" + s.server + ":" + s.pageName;
        s.campaign = "";

        /* Conversion Variables */
        s.eVar1 = "anonymous";
        s.eVar5 = s.channel;
        s.eVar10 = s.prop10;
        s.eVar11 = s.prop11;
        s.eVar17 = "";
        s.eVar23 = s.pageName;
        s.eVar24 = "";
        s.eVar28 = s.prop4;
        s.eVar29 = s.prop9;
        s.eVar46 = s.prop28;

        var s_code = s.t();
        if (s_code) document.write(s_code);
    </script>

            <script src="/Scripts/homeTecoloco.js"></script>






            <div id="updateCandidateData">

            </div>
            
    <script>
                    $('.document').ready(
                        function () {
                            showSearchIconOnScroll(".phone-btnSearch-sub2", 130);
                        }
                    )
    </script>


        </div>

        
        
        <script src="/Scripts/popups-responsive.js" type="text/javascript"></script>
        <script src="/Scripts/2016/jquery.cookie.js" type="text/javascript"></script>
        <script src="/Scripts/2016/videoIniciativa2016.js" type="text/javascript"></script>

 

        <div>
            <a class="b-close"><i class="fa fa-times-circle fa-3x" aria-hidden="true"></i></a>
        </div>

        <div class="hidden-phone">
            <a class="b-close"><i class="fa fa-times-circle fa-3x" aria-hidden="true"></i></a>
        </div>
        
        <div class="overlay hidden-phone">
            <div class="modal-video">
                <div class="video-wrapper">

                </div>
            </div>
            <div class="close-video">

                <i class="fa fa-times fa-lg" aria-hidden="true"></i>

            </div>
        </div>   

        <div class="responsive-ads hidden-desktop ">

            <div class="container">

                <h2>Descarga nuestra app, disponible en:</h2>

                <ul>

                    <li class="pull-left"><a href="https://itunes.apple.com/us/app/tecoloco.com-bolsa-trabajo/id1134960846" target="_blank"><img src="/Content/images/appStore.png" alt="App Store"></a></li>
                    <li class="pull-left"><a href="https://play.google.com/store/apps/details?id=com.stepstone.tecoloco&amp;hl=es" target="_blank"><img src="/Content/images/googlePlay.png" alt="App Store"></a></li>

                </ul>
                <a class="b-close cerrarResponsiveAd"><i class="fa fa-times-circle" aria-hidden="true"></i></a>
            </div>

        </div>




       

        <script>

            /*Llamado de URL videos*/

            $('document').ready(
    function(){



        onClickShowVideo('#btnVideoTrigger2', 'uAW1Fg0JY60?rel=0&autoplay=1', '.video-wrapper');

        onClickShowVideo('#btnVideoTrigger', 'h10qBgyXDn4?rel=0&autoplay=1', '.video-wrapper');

        onClickCloseVideo('.close-video');



    }
);

        </script>

    </body>
</html>