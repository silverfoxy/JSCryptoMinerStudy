<!DOCTYPE html PUBLIC "-//W3C//DTD HTML+RDFa 1.1//EN">
<html lang="es" dir="ltr" version="HTML+RDFa 1.1"
  xmlns:content="http://purl.org/rss/1.0/modules/content/"
  xmlns:dc="http://purl.org/dc/terms/"
  xmlns:foaf="http://xmlns.com/foaf/0.1/"
  xmlns:og="http://ogp.me/ns#"
  xmlns:rdfs="http://www.w3.org/2000/01/rdf-schema#"
  xmlns:sioc="http://rdfs.org/sioc/ns#"
  xmlns:sioct="http://rdfs.org/sioc/types#"
  xmlns:skos="http://www.w3.org/2004/02/skos/core#"
  xmlns:xsd="http://www.w3.org/2001/XMLSchema#">
<head profile="http://www.w3.org/1999/xhtml/vocab">
  <meta http-equiv="Content-Type" content="text/html; charset=utf-8" />
<link rel="shortcut icon" href="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/fav.png" type="image/png" />
<meta name="viewport" content="width=device-width, initial-scale=1, maximum-scale=1, minimum-scale=1, user-scalable=yes" />
<meta name="description" content="Conectate con nuestros planes pospago y prepago para celulares, Internet móvil con la mejor Red LTE 4G de todo El Salvador y las mejores promociones que Tigo tiene para vos. Solo debés Ingresar aquí para conocer ¡todo un mundo digital que espera por ti!" />
<meta name="generator" content="Drupal 7 (http://drupal.org)" />
<link rel="canonical" href="https://www.tigo.com.sv" />
<link rel="shortlink" href="https://www.tigo.com.sv/" />
  <title>Tigo El Salvador | Planes Pospago, Prepago e Internet Móvil</title>
  <style type="text/css" media="all">
@import url("https://www.tigo.com.sv/modules/system/system.base.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/system/system.menus.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/system/system.messages.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/system/system.theme.css?p5wf0x");
</style>
<style type="text/css" media="all">
@import url("https://www.tigo.com.sv/modules/field/theme/field.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/node/node.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/picture/picture_wysiwyg.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/search/search.css?p5wf0x");
@import url("https://www.tigo.com.sv/modules/user/user.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/views/css/views.css?p5wf0x");
</style>
<style type="text/css" media="all">
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/ctools/css/ctools.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/messageclose/css/messageclose.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_dynamic_background/css/tigosmart_dynamic_background.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/tigowebcorp.sv/files/css/social_icons.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/tigowebcorp.sv/files/tigo_graphic_menu_icons/tigo_graphic_menu_icons.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_custom_pages/plugins/layouts/onecol/onecol.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/field_group/field_group.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/field_collection/field_collection.theme.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/flexslider/assets/css/flexslider_img.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/libraries/flexslider/flexslider.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/fonts/font-awesome/css/font-awesome.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/css/bootstrap.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/css/base.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/css/default.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/css/compatibility.css?p5wf0x");
</style>
<style type="text/css" media="all">
@import url("https://www.tigo.com.sv/sites/all/modules/custom/tigo_graphic_menu/css/tigo_menu_themes.css?p5wf0x");
</style>
<style type="text/css" media="all">
@import url("https://www.tigo.com.sv/sites/all/themes/omega/alpha/css/alpha-reset.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/alpha/css/alpha-mobile.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/alpha/css/alpha-alpha.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/formalize.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/omega-text.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/omega-branding.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/omega-menu.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/omega-forms.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/omega/css/omega-visuals.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/global.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/moni.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/style.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/tigowebcorp.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/tigowebcorp.sv.css?p5wf0x");
</style>

<!--[if (lt IE 9)&(!IEMobile)]>
<style type="text/css" media="all">
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/tigo-smart-alpha-default.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/alpha/css/grid/alpha_default/fluid/alpha-default-fluid-12.css?p5wf0x");
</style>
<![endif]-->

<!--[if gte IE 9]><!-->
<style type="text/css" media="all and (min-width: 980px) and (min-device-width: 980px), all and (max-device-width: 1024px) and (min-width: 1024px) and (orientation:landscape)">
@import url("https://www.tigo.com.sv/sites/all/themes/tigo_smart/css/tigo-smart-alpha-default.css?p5wf0x");
@import url("https://www.tigo.com.sv/sites/all/themes/omega/alpha/css/grid/alpha_default/fluid/alpha-default-fluid-12.css?p5wf0x");
</style>
<!--<![endif]-->
  <script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/jquery_update/replace/jquery/1.7/jquery.min.js?v=1.7.2"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/misc/drupal.js?p5wf0x"></script>
<script type="text/javascript">
<!--//--><![CDATA[//><!--
document.createElement( "picture" );
//--><!]]>
</script>
<script type="text/javascript">
<!--//--><![CDATA[//><!--
delete Drupal.behaviors.tbMegaMenuAction
//--><!]]>
</script>
<script type="text/javascript">
<!--//--><![CDATA[//><!--
jQuery.extend(Drupal.settings, {"basePath":"\/","pathPrefix":"","ajaxPageState":{"theme":"tigo_smart","theme_token":"-Q91lr1elfABjHqIhnzXR5BdSWKbDa6vM16ifT_w3YA","js":{"sites\/all\/libraries\/respondjs\/respond.min.js":1,"misc\/jquery.once.js":1,"sites\/all\/modules\/contrib\/jquery_update\/replace\/ui\/ui\/minified\/jquery.ui.effect.min.js":1,"sites\/all\/modules\/contrib\/jquery_update\/replace\/ui\/ui\/minified\/jquery.ui.effect-slide.min.js":1,"sites\/all\/modules\/contrib\/picture\/picturefill2\/picturefill.min.js":1,"sites\/all\/modules\/contrib\/picture\/picture.min.js":1,"sites\/all\/modules\/custom\/tigo_graphic_menu\/js\/tigo_menu_themes.js":1,"sites\/all\/modules\/contrib\/messageclose\/js\/messageclose.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/detectmobilebrowser.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/jquery.wait.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/jquery.fittext.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/tigosmart_customjs.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/tigosmart_js.js":1,"sites\/all\/modules\/custom\/tigosmart_customjs\/waypoints.min.js":1,"sites\/all\/modules\/custom\/tigosmart_custom_pages\/js\/panel_ajax_loader.js":1,"sites\/all\/modules\/contrib\/field_group\/field_group.js":1,"sites\/all\/libraries\/flexslider\/jquery.flexslider-min.js":1,"sites\/all\/modules\/contrib\/flexslider\/assets\/js\/flexslider.load.js":1,"sites\/all\/modules\/contrib\/tb_megamenu\/js\/tb-megamenu-frontend.js":1,"sites\/all\/modules\/custom\/features\/display_data_set_lists_fragment\/js\/display_data_set_lists_fragment.js":1,"sites\/all\/modules\/contrib\/tb_megamenu\/js\/tb-megamenu-touch.js":1,"sites\/all\/themes\/omega\/omega\/js\/jquery.formalize.js":1,"sites\/all\/themes\/omega\/omega\/js\/omega-mediaqueries.js":1,"sites\/all\/themes\/tigo_smart\/js\/jquery.mmenu.js":1,"sites\/all\/themes\/tigo_smart\/js\/tigowebcorp.scripts.js":1,"sites\/all\/modules\/contrib\/jquery_update\/replace\/jquery\/1.7\/jquery.min.js":1,"misc\/drupal.js":1,"0":1,"1":1},"css":{"modules\/system\/system.base.css":1,"modules\/system\/system.menus.css":1,"modules\/system\/system.messages.css":1,"modules\/system\/system.theme.css":1,"modules\/field\/theme\/field.css":1,"modules\/node\/node.css":1,"sites\/all\/modules\/contrib\/picture\/picture_wysiwyg.css":1,"modules\/search\/search.css":1,"modules\/user\/user.css":1,"sites\/all\/modules\/contrib\/views\/css\/views.css":1,"sites\/all\/modules\/contrib\/ctools\/css\/ctools.css":1,"sites\/all\/modules\/contrib\/messageclose\/css\/messageclose.css":1,"sites\/all\/modules\/custom\/tigosmart_dynamic_background\/css\/tigosmart_dynamic_background.css":1,"public:\/\/css\/social_icons.css":1,"public:\/\/tigo_graphic_menu_icons\/tigo_graphic_menu_icons.css":1,"sites\/all\/modules\/custom\/tigosmart_custom_pages\/plugins\/layouts\/onecol\/onecol.css":1,"sites\/all\/modules\/contrib\/field_group\/field_group.css":1,"sites\/all\/modules\/contrib\/field_collection\/field_collection.theme.css":1,"sites\/all\/modules\/contrib\/flexslider\/assets\/css\/flexslider_img.css":1,"sites\/all\/libraries\/flexslider\/flexslider.css":1,"sites\/all\/modules\/contrib\/tb_megamenu\/fonts\/font-awesome\/css\/font-awesome.css":1,"sites\/all\/modules\/contrib\/tb_megamenu\/css\/bootstrap.css":1,"sites\/all\/modules\/contrib\/tb_megamenu\/css\/base.css":1,"sites\/all\/modules\/contrib\/tb_megamenu\/css\/default.css":1,"sites\/all\/modules\/contrib\/tb_megamenu\/css\/compatibility.css":1,"sites\/all\/modules\/custom\/tigo_graphic_menu\/css\/tigo_menu_themes.css":1,"sites\/all\/themes\/omega\/alpha\/css\/alpha-reset.css":1,"sites\/all\/themes\/omega\/alpha\/css\/alpha-mobile.css":1,"sites\/all\/themes\/omega\/alpha\/css\/alpha-alpha.css":1,"sites\/all\/themes\/omega\/omega\/css\/formalize.css":1,"sites\/all\/themes\/omega\/omega\/css\/omega-text.css":1,"sites\/all\/themes\/omega\/omega\/css\/omega-branding.css":1,"sites\/all\/themes\/omega\/omega\/css\/omega-menu.css":1,"sites\/all\/themes\/omega\/omega\/css\/omega-forms.css":1,"sites\/all\/themes\/omega\/omega\/css\/omega-visuals.css":1,"sites\/all\/themes\/tigo_smart\/css\/global.css":1,"sites\/all\/themes\/tigo_smart\/css\/moni.css":1,"sites\/all\/themes\/tigo_smart\/css\/style.css":1,"sites\/all\/themes\/tigo_smart\/css\/tigowebcorp.css":1,"sites\/all\/themes\/tigo_smart\/css\/tigowebcorp.sv.css":1,"ie::fluid::sites\/all\/themes\/tigo_smart\/css\/tigo-smart-alpha-default.css":1,"ie::fluid::sites\/all\/themes\/omega\/alpha\/css\/grid\/alpha_default\/fluid\/alpha-default-fluid-12.css":1,"fluid::sites\/all\/themes\/tigo_smart\/css\/tigo-smart-alpha-default.css":1,"sites\/all\/themes\/omega\/alpha\/css\/grid\/alpha_default\/fluid\/alpha-default-fluid-12.css":1}},"tigosmart_custom_pages_ajax_panel":{"cid":"tigosmart_cp_panel_ajax:panel_context:page-pagina_principal::page_pagina_principal_panel_context::::","width_mobile":767},"field_group":{"div":"desktop"},"flexslider":{"optionsets":{"default":{"namespace":"flex-","selector":".slides \u003E li","easing":"swing","direction":"horizontal","reverse":false,"smoothHeight":false,"startAt":0,"animationSpeed":600,"initDelay":0,"useCSS":true,"touch":true,"video":false,"keyboard":true,"multipleKeyboard":false,"mousewheel":false,"controlsContainer":".flex-control-nav-container","sync":"","asNavFor":"","itemWidth":0,"itemMargin":0,"minItems":0,"maxItems":0,"move":0,"animation":"fade","slideshow":true,"slideshowSpeed":7000,"directionNav":true,"controlNav":true,"prevText":"Previous","nextText":"Next","pausePlay":false,"pauseText":"Pause","playText":"Play","randomize":false,"thumbCaptions":false,"thumbCaptionsBoth":false,"animationLoop":true,"pauseOnAction":true,"pauseOnHover":false,"manualControls":""}},"instances":{"flexslider-1":"default"}},"data_set_lists":[{"url":"http:\/\/www.tigobusiness.com.sv\/","el":"content-setlists-theme-vertical-blue-bg-with-btn-50","class_name":"content-setlists-theme-vertical-blue-bg-with-btn-entire-clickable"},{"url":"http:\/\/internet.tigo.com.sv","el":"content-setlists-theme-vertical-blue-bg-with-btn-52","class_name":"content-setlists-theme-vertical-blue-bg-with-btn-entire-clickable"},{"url":"https:\/\/www.tigo.com.sv\/tigo\/postpago","el":"content-setlists-theme-vertical-blue-bg-with-btn-53","class_name":"content-setlists-theme-vertical-blue-bg-with-btn-entire-clickable"},{"url":"http:\/\/www.tigomoney.com.sv\/","el":"content-setlists-theme-2cols-transparent-bg-stt-link-54","class_name":"content-setlists-theme-2cols-transparent-bg-stt-link-entire-clickable"},{"url":"https:\/\/www.tigo.com.sv\/renova-tu-plan","el":"content-setlists-theme-2cols-transparent-bg-stt-link-55","class_name":"content-setlists-theme-2cols-transparent-bg-stt-link-entire-clickable"},{"url":"https:\/\/www.tigo.com.sv\/portabilidad","el":"content-setlists-theme-2cols-transparent-bg-stt-link-56","class_name":"content-setlists-theme-2cols-transparent-bg-stt-link-entire-clickable"}],"omega":{"layouts":{"primary":"fluid","order":["fluid"],"queries":{"fluid":"all and (min-width: 980px) and (min-device-width: 980px), all and (max-device-width: 1024px) and (min-width: 1024px) and (orientation:landscape)"}}}});
//--><!]]>
</script>
  <!--[if lt IE 9]><script src="http://html5shiv.googlecode.com/svn/trunk/html5.js"></script><![endif]-->
</head>
<body class="html front not-logged-in page-home tigosmart-custom-body-class dl-class dd-desktop device-detected" id="dark-blue">
<!-- Google Tag Manager -->
<noscript><iframe src="//www.googletagmanager.com/ns.html?id=GTM-W3PB5W" height="0" width="0" style="display:none;visibility:hidden"></iframe></noscript>
<script type="text/javascript">(function(w,d,s,l,i){w[l]=w[l]||[];w[l].push({'gtm.start':new Date().getTime(),event:'gtm.js'});var f=d.getElementsByTagName(s)[0];var j=d.createElement(s);var dl=l!='dataLayer'?'&l='+l:'';j.src='//www.googletagmanager.com/gtm.js?id='+i+dl;j.type='text/javascript';j.async=true;f.parentNode.insertBefore(j,f);})(window,document,'script','dataLayer','GTM-W3PB5W');</script>
<!-- End Google Tag Manager -->
    <div id="skip-link">
    <a href="#main-content" class="element-invisible element-focusable">saltar el contenido principal </a>
  </div>
    <div class="page clearfix" id="page">
      <header id="section-header" class="section section-header">
  <div id="zone-user-wrapper" class="zone-wrapper zone-user-wrapper clearfix">  
  <div id="zone-user" class="zone zone-user clearfix container-12">
    <div class="grid-12 region region-user-first" id="region-user-first">
  <div class="region-inner region-user-first-inner">
    <div class="block block-menu top-menu block-menu-tigosmart-top-menu block-menu-menu-tigosmart-top-menu odd block-without-title" id="block-menu-menu-tigosmart-top-menu">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <ul class="menu"><li class="first leaf active-trail"><a href="/" class="active-trail active">Móvil</a></li>
<li class="leaf"><a href="http://www.tigostar.com.sv/"> Residencial </a></li>
<li class="leaf"><a href="http://www.tigobusiness.com.sv/">Tigo Business</a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/tigo-money-0">Tigo Money</a></li>
<li class="leaf"><a href="http://www.tigomusic.sv/" class="tigo-productos-link">TIGO MUSIC</a></li>
<li class="last leaf"><a href="https://www.tigo.com.sv/tigosports" class="tigo-productos-link">TIGO SPORTS</a></li>
</ul>    </div>
  </div>
</div><div class="block block-tb-megamenu block-user-menu block-tb-megamenu-user-menu even block-without-title" id="block-tb-megamenu-user-menu">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div  class="tb-megamenu tb-megamenu-user-menu tb-megamenu-main-menu" class="tb-megamenu tb-megamenu-user-menu tb-megamenu-main-menu">
      <button data-target=".nav-collapse" data-toggle="collapse" class="btn btn-navbar tb-megamenu-button" type="button">
      <i class="icon-reorder"></i>
    </button>
    <div class="nav-collapse collapse always-show">
    <div class="div-dropdown-toggle left"></div>
<ul  class="tb-megamenu-nav nav level-0 items-4" class="tb-megamenu-nav nav level-0 items-4">
  <li  data-id="1353" data-level="1" data-type="menu_item" data-class="" data-xicon="" data-caption="" data-alignsub="" data-group="0" data-hidewcol="0" data-hidesub="0" class="tb-megamenu-item level-1 mega" class="tb-megamenu-item level-1 mega">
    <a href="https://compras.tigo.com.sv/" class="tienda-online">
        Tienda Online          </a>
  </li>

<li  data-id="1626" data-level="1" data-type="menu_item" data-class="" data-xicon="" data-caption="" data-alignsub="" data-group="0" data-hidewcol="0" data-hidesub="0" class="tb-megamenu-item level-1 mega" class="tb-megamenu-item level-1 mega">
    <a href="https://ayuda.tigo.com.sv/hc/es/" class="">
        Atención al Cliente          </a>
  </li>

<li  data-id="1883" data-level="1" data-type="menu_item" data-class="" data-xicon="" data-caption="" data-alignsub="" data-group="0" data-hidewcol="0" data-hidesub="0" class="tb-megamenu-item level-1 mega" class="tb-megamenu-item level-1 mega">
    <a href="http://micuenta.tigo.com.sv/" class="">
        Mi Cuenta          </a>
  </li>
</ul>
<div class="div-dropdown-toggle right"></div>
      </div>
  </div>
    </div>
  </div>
</div>  </div>
</div>  </div>
</div><div id="zone-header-wrapper" class="zone-wrapper zone-header-wrapper clearfix">  
  <div id="zone-header" class="zone zone-header clearfix container-12">
    <div class="page-mask">
      <div class="page-loader">
      </div>
</div>
<!-- Page Mask End _Finalizar loader de la pagina_ -->
  <div id="navmobile" >
    <div class="mm-menu-content">
    <div class="block block-menu main-menu-mobile block- block-menu-main-menu-mobile block-menu-menu-main-menu-mobile odd block-without-title" id="block-menu-menu-main-menu-mobile">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <ul class="menu"><li class="first leaf active-trail"><a href="/" class="active-trail active">Inicio</a></li>
<li class="leaf"><a href="/tigo/postpago">Pospago</a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/tigo/prepago">Prepago</a></li>
<li class="leaf"><a href="http://internet.tigo.com.sv/">Paquetigos</a></li>
<li class="leaf"><a href="/tigo/telefonos">Smartphones</a></li>
<li class="expanded has-submenu"><a href="javascript: void(0);">Apps y Servicios</a><ul class="menu"><li class="first leaf"><a href="/mi-tigo-app">Mi Tigo</a></li>
<li class="leaf"><a href="/shop">Tigo Shop</a></li>
<li class="leaf"><a href="/smart-apps">Smartapps</a></li>
<li class="leaf"><a href="http://deezer.tigo.com.bo/">Tigo Music</a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/tigosports">Tigo Sports</a></li>
<li class="last leaf"><a href="/tigo-money-0">Tigo Money</a></li>
</ul></li>
<li class="leaf"><a href="https://compras.tigo.com.sv/" class="tienda-online">Tienda Online</a></li>
<li class="leaf"><a href="https://ayuda.tigo.com.sv/hc/es/">Ayuda</a></li>
<li class="leaf"><a href="http://micuenta.tigo.com.sv/">Mi Cuenta</a></li>
<li class="last expanded has-submenu"><a href="#">Otros Productos Tigo</a><ul class="menu"><li class="first last leaf"><a href="http://www.tigostar.com.sv/">Tigo Star</a></li>
</ul></li>
</ul>    </div>
  </div>
</div><div class="block block-block block- block-4 block-block-4 even block-without-title" id="block-block-4">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <script>
<!--//--><![CDATA[// ><!--


jQuery(function ($) {
 
  $("ul li.leaf a div").css({'font-family':'Roboto, sans-serif', 'font-size': '15px', 'color': '#fff', 'padding':'0'});

});

//--><!]]>
</script>    </div>
  </div>
</div>    </div>
  </div>
<div class="grid-12 region region-header-logo" id="region-header-logo">
  <div class="region-inner region-header-logo-inner">
    <div class="block block-block header-mobile block-3 block-block-3 odd block-without-title" id="block-block-3">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="mobile-btn-wrapper"><a id="mobile-menu-btn" href="#navmobile">MENU</a></div>
<div id="logo-mobile"><a href="/"><img src="/sites/tigowebcorp.bo/files/logo.svg" /></a></div>
    </div>
  </div>
</div><div class="block block-delta-blocks block-logo block-delta-blocks-logo even block-without-title" id="block-delta-blocks-logo">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="logo-img"><a href="/" id="logo" title="Return to the Movil Web home page"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/logo.svg" alt="Movil Web" /></a></div>    </div>
  </div>
</div><div class="block block-menu block-menu-menu-header-logo block-menu-menu-menu-header-logo odd block-without-title" id="block-menu-menu-menu-header-logo">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <ul class="menu menu-theme-icons-desktop"><li class="first leaf"><a href="/tigo/postpago">Pospago</a></li>
<li class="leaf"><a href="/Tigo/prepago"><div class='tigo-graphic-menu-icons-1699 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Prepago</div></a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/shop"><div class='tigo-graphic-menu-icons-1700 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Paquetigos</div></a></li>
<li class="leaf"><a href="/tigo/telefonos"><div class='tigo-graphic-menu-icons-1701 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Smartphones</div></a></li>
<li class="last expanded has-submenu"><a href="javascript: void(0);">Apps y Servicios</a><ul class="menu"><li class="first leaf"><a href="/mi-tigo-app"><div class='tigo-graphic-menu-icons-1703 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Mi Tigo</div><div class='caption-menu-theme-icons-desktop'>Consulta tu saldo disponible y el consumo de tus servicios desde tu smartphone.</div></a></li>
<li class="leaf"><a href="/shop"><div class='tigo-graphic-menu-icons-1704 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Tigo Shop</div><div class='caption-menu-theme-icons-desktop'>Compra Paquetigos para tu smartphone de manera fácil, rápida y segura.</div></a></li>
<li class="leaf"><a href="/smart-apps"><div class='tigo-graphic-menu-icons-2068 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Smartapps</div><div class='caption-menu-theme-icons-desktop'>Compra Paquetigos para tu smartphone de manera fácil, rápida y segura.</div></a></li>
<li class="leaf"><a href="http://www.tigomusic.sv "><div class='tigo-graphic-menu-icons-1977 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Tigo Music</div><div class='caption-menu-theme-icons-desktop'>Enterate las últimas noticias del mundo de la música y escuchá las mejores playlists.</div></a></li>
<li class="leaf"><a href="https://wwwold.tigo.com.sv/tigosports"><div class='tigo-graphic-menu-icons-2069 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Tigo Sports</div><div class='caption-menu-theme-icons-desktop'>Todas las noticias del deporte y las mejores repeticiones en un solo lugar.</div></a></li>
<li class="last leaf"><a href="http://www.tigomoney.com.sv/"><div class='tigo-graphic-menu-icons-2071 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-desktop'>Tigo Money</div><div class='caption-menu-theme-icons-desktop'>Controla tu billetera digital, realiza pagos de servicios y recarga tu saldo.</div></a></li>
</ul></li>
</ul>    </div>
  </div>
</div>  </div>
</div>  </div>
</div></header>    
      <section id="section-content" class="section section-content">
  <div id="zone-content-wrapper" class="zone-wrapper zone-content-wrapper clearfix">  
  <div id="zone-content" class="zone zone-content clearfix container-12">    
        
        <div class="grid-12 region region-content" id="region-content">
  <div class="region-inner region-content-inner">
    <a id="main-content"></a>
                        <div class="block block-system block-main block-system-main odd block-without-title" id="block-system-main">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class='tigosmart-custom-page-content'><div class="panel-display panel-1col clearfix" >
  <div class="panel-panel panel-col">
    <div><div class="block block-bean block-banner-11082017 block-bean-banner-11082017 odd block-without-title slideshow_multi_line_banner slideshow-multi-line-banner-block-bean" id="block-bean-banner-11082017">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="entity entity-bean bean-slideshow-multi-line-banner clearfix" about="/block/banner-11082017" typeof="" class="entity entity-bean bean-slideshow-multi-line-banner">

  <div class="content">
    <h2 class="bean-title"></h2>
<div  id="flexslider-1" class="flexslider">
  <ul class="slides"><li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/330" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/330"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/plan-recarga-mensual"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/BannersWeb-PospTigo-OM_0.png" width="1280" height="375" alt="Recarga mensual Tigo" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-330 multi-line-banner-box-float-left multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-left</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/290" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/290"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="http://www.tigostar.com.sv/entretenimientotigo"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/TSV_B2S_HOME_DESKT_0.jpg" width="1280" height="375" alt="Tv Digital para Vivir el Cine en tu Casa " /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-290 multi-line-banner-box-float-left multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-left</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/321" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/321"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/samsung-galaxy-s9"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/samsung-galaxy-s9-banner-desk_0_0.jpg" width="1280" height="375" alt="Smartphone Samsung Galaxy S9" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-321 multi-line-banner-box-float-left multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-left</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/300" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/300"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/ofertas_pospago"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/TSV_ECOMMERCE_HOMEDESK_SJ2.jpg" width="1280" height="375" alt="Promoción del Smartphone Samsung J2 Prime" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-300 multi-line-banner-box-float-left multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-left</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/251" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/251"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/ofertas_pospago"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/TSV_ECOMMERCE_HOMEDESK_LGK8.jpg" width="1280" height="375" alt="Empieza el Verano con un Smartphone Nuevo en la Red 4G LTE" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-251 multi-line-banner-box-float-bottomleft multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-bottomleft</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/279" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/279"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/ofertas_pospago"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/TSV_ECOMMERCE_HOMEDESK_LGK10.jpg" width="1280" height="375" alt="Empieza el Verano con un Smartphone LG K10 Nuevo" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-279 multi-line-banner-box-float-right multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-right</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
<li><div class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner clearfix" about="/elements_of_fragments/multi_line_banner/257" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-multi-line-banner">

      <h2>
              <a href="/elements_of_fragments/multi_line_banner/257"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-multi-line-banner-bg field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><a href="http://micuenta.tigo.com.sv"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/banner_factura_DESKTOP_0.png" width="1280" height="375" alt="Consulta la Factura de tu Celular Pospago e Internet Móvil" /></a></div></div></div><div class="group-multi-line-banner-wrapper group-multi-line-banner-wrapper-257 multi-line-banner-box-float-right multi-line-banner-box-transparent-bg"><div class="field-collection-container clearfix"><div class="field field-name-field-multi-line-banner-content field-type-field-collection field-label-hidden"><div class="field-items"></div></div></div><div class="field field-name-field-multi-line-banner-box field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-float-right</div></div></div><div class="field field-name-field-multi-line-banner-box-bg field-type-list-text field-label-hidden multi-line-banner-hidden"><div class="field-items"><div class="field-item even">multi-line-banner-box-transparent-bg</div></div></div></div>  </div>
</div>
</li>
</ul></div>
  </div>
</div>
    </div>
  </div>
</div><div class="panel-separator"></div><div class="block block-bean block-destacado28dic block-bean-destacado28dic even block-without-title display_data_setlists display-data-setlists-block-bean" id="block-bean-destacado28dic">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="entity entity-bean bean-display-data-setlists display-data-setlists clearfix" about="/block/destacado28dic" typeof="" class="entity entity-bean bean-display-data-setlists">

  <div class="content">
    <div class="field field-name-field-content-setlists-elements field-type-entityreference field-label-hidden"><div class="field-items"><div class="field-item even"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-vertical-blue-bg content-setlists-theme-vertical-blue-bg-with-btn-50 content-setlists-theme-vertical-blue-bg-stt-no-link clearfix" about="/elements_of_fragments/content_setlists/50" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/50"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-vertical-blue-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/1.%20Boton_B2B%20DESKTOP.png" width="104" height="31" alt="" /></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden"><div class="field-items"><div class="field-item even"><p><strong> Una solución</strong><br />
para tu negocio</p>
</div></div></div><div class="field field-name-field-content-setlists-btn-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="http://www.tigobusiness.com.sv/">CONOCE MÁS</a></div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div><div class="field-item odd"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-vertical-blue-bg content-setlists-theme-vertical-blue-bg-with-btn-52 content-setlists-theme-vertical-blue-bg-stt-no-link clearfix" about="/elements_of_fragments/content_setlists/52" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/52"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-vertical-blue-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/2%20Boton_paquetigo%20DESKTOP.png" width="104" height="31" alt="" /></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden wysiwyg-content"><div class="field-items"><div class="field-item even"><p>Comprá tu paquete <br /><strong>Prepago</strong></p>
</div></div></div><div class="field field-name-field-content-setlists-btn-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="http://internet.tigo.com.sv">COMPRAR</a></div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div><div class="field-item even"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-vertical-blue-bg content-setlists-theme-vertical-blue-bg-with-btn-53 content-setlists-theme-vertical-blue-bg-stt-no-link clearfix" about="/elements_of_fragments/content_setlists/53" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/53"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-vertical-blue-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/3.Boton_pospago%20DESKTOP.png" width="104" height="31" alt="" /></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden wysiwyg-content"><div class="field-items"><div class="field-item even"><p>Ahorrá con tu <br /><strong>plan Pospago</strong></p>
</div></div></div><div class="field field-name-field-content-setlists-btn-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/tigo/postpago">PLANES TIGO</a></div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div></div></div>  </div>
</div>
    </div>
  </div>
</div><div class="panel-separator"></div><div class="block block-bean block-icono28dic block-bean-icono28dic odd block-without-title display_data_setlists display-data-setlists-block-bean" id="block-bean-icono28dic">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="entity entity-bean bean-display-data-setlists display-data-setlists clearfix" about="/block/icono28dic" typeof="" class="entity entity-bean bean-display-data-setlists">

  <div class="content">
    <div class="field field-name-field-content-setlists-elements field-type-entityreference field-label-hidden"><div class="field-items"><div class="field-item even"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-2cols-transparent-bg content-setlists-theme-2cols-transparent-bg-without-btn content-setlists-theme-2cols-transparent-bg-stt-link-54 clearfix" about="/elements_of_fragments/content_setlists/54" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/54"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-2cols-transparent-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/Tigo%20Money%20-%20Desktop.png" width="48" height="61" alt="" /></div></div></div><div class="field field-name-field-content-setlists-stt-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="http://www.tigomoney.com.sv/">Tigo Money</a></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden wysiwyg-content"><div class="field-items"><div class="field-item even"><p>Tu billetera electrónica<br />
desde tu smartphone </p>
</div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">1</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div><div class="field-item odd"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-2cols-transparent-bg content-setlists-theme-2cols-transparent-bg-without-btn content-setlists-theme-2cols-transparent-bg-stt-link-55 clearfix" about="/elements_of_fragments/content_setlists/55" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/55"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-2cols-transparent-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/renova-planV2.png" width="48" height="61" alt="" /></div></div></div><div class="field field-name-field-content-setlists-stt-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/renova-tu-plan">Renová tu Plan</a></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden"><div class="field-items"><div class="field-item even"><p>Seguí disfrutando todos tus beneficios pospago <a href="https://www.tigo.com.sv/renova-tu-plan">Aquí</a></p>
</div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">1</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div><div class="field-item even"><div class="entity entity-elements-of-fragments elements-of-fragments-content-setlists content-setlists-theme-2cols-transparent-bg content-setlists-theme-2cols-transparent-bg-without-btn content-setlists-theme-2cols-transparent-bg-stt-link-56 clearfix" about="/elements_of_fragments/content_setlists/56" typeof="" class="entity entity-elements-of-fragments elements-of-fragments-content-setlists">

      <h2>
              <a href="/elements_of_fragments/content_setlists/56"></a>
          </h2>
  
  <div class="content">
    <div class="field field-name-field-content-setlists-theme field-type-list-text field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">content-setlists-theme-2cols-transparent-bg</div></div></div><div class="field field-name-field-content-setlists-image-img field-type-image field-label-hidden"><div class="field-items"><div class="field-item even"><img typeof="foaf:Image" src="https://www.tigo.com.sv/sites/tigowebcorp.sv/files/Portabilidad-Desktop.png" width="48" height="61" alt="" /></div></div></div><div class="field field-name-field-content-setlists-stt-link field-type-link-field field-label-hidden"><div class="field-items"><div class="field-item even"><a href="https://www.tigo.com.sv/portabilidad">Portabilidad</a></div></div></div><div class="field field-name-field-content-setlists-desc-txt field-type-text-long field-label-hidden"><div class="field-items"><div class="field-item even"><p>Pasate ya al mejor internet LTE 4G</p>
</div></div></div><div class="field field-name-field-content-setlists-sttl-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">1</div></div></div><div class="field field-name-field-content-setlists-head-depe field-type-list-boolean field-label-hidden content-setlists-hidden"><div class="field-items"><div class="field-item even">0</div></div></div>  </div>
</div>
</div></div></div>  </div>
</div>
    </div>
  </div>
</div></div>
  </div>
</div>
</div>    </div>
  </div>
</div>      </div>
</div>  </div>
</div><div id="zone-content-bottom-wrapper" class="zone-wrapper zone-content-bottom-wrapper clearfix">  
  <div id="zone-content-bottom" class="zone zone-content-bottom clearfix container-12">
    <div class="grid-12 region region-content-bottom-first" id="region-content-bottom-first">
  <div class="region-inner region-content-bottom-first-inner">
    <div class="block block-menu otros-productos-menu block-menu-otros-productos-mobile block-menu-menu-otros-productos-mobile odd block-without-title" id="block-menu-menu-otros-productos-mobile">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <ul class="menu"><li class="first last expanded has-submenu"><a href="javascript: void(0);">Otros Productos</a><ul class="menu"><li class="first leaf"><a href="/tigo">TIGO</a></li>
<li class="leaf"><a href="http://www.tigostar.com.sv/"> RESIDENCIAL</a></li>
<li class="leaf"><a href="http://tigobusiness.com.sv/">TIGO BUSINESS</a></li>
<li class="leaf"><a href="http://www.tigomoney.com.sv/">TIGO MONEY</a></li>
<li class="leaf"><a href="http://www.tigomusic.sv/">TIGO MUSIC</a></li>
<li class="last leaf"><a href="http://www.tigo.com.sv/tigosports">TIGO SPORTS</a></li>
</ul></li>
</ul>    </div>
  </div>
</div>  </div>
</div>  </div>
</div></section>    
  
      <footer id="section-footer" class="section section-footer">
  <div id="zone-footer-blocks-wrapper" class="zone-wrapper zone-footer-blocks-wrapper clearfix">  
  <div id="zone-footer-blocks" class="zone zone-footer-blocks clearfix container-12">
    <div class="grid-3 region region-footer-first" id="region-footer-first">
  <div class="region-inner region-footer-first-inner">
    <section class="block block-menu block-menu-un-estilo-de-vida-digital block-menu-menu-un-estilo-de-vida-digital odd" id="block-menu-menu-un-estilo-de-vida-digital">
  <div class="block-inner clearfix">
              <h2 class="block-title">Mundo Tigo </h2>
            
    <div class="content clearfix">
      <ul class="menu menu-theme-icons-mobile"><li class="first leaf"><a href="https://www.tigo.com.sv/tigo-corporativo"><div class='tigo-graphic-menu-icons-1628 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-mobile'>Historia Corporativa</div></a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/content/responsabilidad-corporativa"><div class='tigo-graphic-menu-icons-1630 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-mobile'>Responsabilidad Social</div></a></li>
<li class="leaf"><a href="http://crianzatecnologica.org/" target="_blank"><div class='tigo-graphic-menu-icons-2465 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-mobile'>Crianza Digital</div></a></li>
<li class="leaf"><a href="/terminos"><div class='tigo-graphic-menu-icons-2519 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-mobile'>Términos y condiciones</div></a></li>
<li class="last leaf"><a href="https://www.tigo.com.sv/promociones-vigentes"><div class='tigo-graphic-menu-icons-0 tigo-graphic-menu-icons'></div><div class='title-menu-theme-icons-mobile'>Promociones Vigentes</div></a></li>
</ul>    </div>
  </div>
</section>  </div>
</div><div class="grid-3 region region-footer-second" id="region-footer-second">
  <div class="region-inner region-footer-second-inner">
    <section class="block block-menu block-menu-apps block-menu-menu-apps odd" id="block-menu-menu-apps">
  <div class="block-inner clearfix">
              <h2 class="block-title">TIGO APPS</h2>
            
    <div class="content clearfix">
      <ul class="menu"><li class="first leaf"><a href="/shop">Tigo Shop</a></li>
<li class="leaf"><a href="/tigo-money-0">Tigo Money </a></li>
<li class="leaf"><a href="/mi-tigo-app">Mi Tigo</a></li>
<li class="leaf"><a href="https://www.tigo.com.sv/tigosports">Tigo Sports </a></li>
<li class="last leaf"><a href="/smart-apps">SmartApps</a></li>
</ul>    </div>
  </div>
</section>  </div>
</div><div class="grid-3 region region-footer-third" id="region-footer-third">
  <div class="region-inner region-footer-third-inner">
    <section class="block block-menu block-menu-atenci-n-al-cliente block-menu-menu-atenci-n-al-cliente odd" id="block-menu-menu-atenci-n-al-cliente">
  <div class="block-inner clearfix">
              <h2 class="block-title">Atención al cliente</h2>
            
    <div class="content clearfix">
      <ul class="menu"><li class="first leaf"><a href="https://ayuda.tigo.com.sv/hc/es/">Preguntas frecuentes </a></li>
<li class="leaf"><a href="https://ayuda.tigo.com.sv/hc/es/requests/new?ticket_form_id=577188">Escribinos</a></li>
<li class="leaf"><a href="https://wwwold.tigo.com.sv/personas/horarios-de-tiendas-tigo">Horarios de tiendas</a></li>
<li class="last leaf"><a href="javascript: void(0);"> *611 Gratis desde tu Tigo</a></li>
</ul>    </div>
  </div>
</section>  </div>
</div>  </div>
</div><div id="zone-footer-wrapper" class="zone-wrapper zone-footer-wrapper clearfix">  
  <div id="zone-footer" class="zone zone-footer clearfix container-12">
    <div class="grid-12 region region-footer-bottom-first" id="region-footer-bottom-first">
  <div class="region-inner region-footer-bottom-first-inner">
    <div class="block block-block block-1 block-block-1 odd block-without-title" id="block-block-1">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <p>Esta empresa está regulada y fiscalizada por la Autoridad de Regulación y Fiscalización de Telecomunicaciones y Transportes.<br />
Tigo Copyright © 2018. Tigo El Salvador. Todos los derechos reservados.</p>
    </div>
  </div>
</div>  </div>
</div><div class="grid-12 region region-footer-bottom-second" id="region-footer-bottom-second">
  <div class="region-inner region-footer-bottom-second-inner">
    <div class="block block-tigosmart-social-networks block-block-tigosmart-social-networks block-tigosmart-social-networks-block-tigosmart-social-networks odd block-without-title" id="block-tigosmart-social-networks-block-tigosmart-social-networks">
  <div class="block-inner clearfix">
                
    <div class="content clearfix">
      <div class="message-header-social-network">Síguenos en:</div>
<ul class="items-social-network" />
<li class="item-social item-social-1"><a href="https://www.facebook.com/tigosv/" target="_blank"><span class="sprite-icon Facebook social-network-Facebook" />
</a></li>
<li class="item-social item-social-2"><a href="https://twitter.com/tigoelsalvador?lang=es" target="_blank"><span class="sprite-icon Twitter  social-network-Twitter-" />
</a></li>
<li class="item-social item-social-3"><a href="https://www.instagram.com/tigoelsalvador/" target="_blank"><span class="sprite-icon Instagram  social-network-Instagram-" />
</a></li>
<li class="item-social item-social-4"><a href="https://www.youtube.com/user/TigoElsalvador" target="_blank"><span class="sprite-icon You Tube social-network-You-Tube" />
</a></li>
    </div>
  </div>
</div>  </div>
</div>  </div>
</div></footer>  </div>  <script type="text/javascript" src="https://www.tigo.com.sv/sites/all/libraries/respondjs/respond.min.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/misc/jquery.once.js?v=1.2"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/jquery_update/replace/ui/ui/minified/jquery.ui.effect.min.js?v=1.10.2"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/jquery_update/replace/ui/ui/minified/jquery.ui.effect-slide.min.js?v=1.10.2"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/picture/picturefill2/picturefill.min.js?v=2.3.1"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/picture/picture.min.js?v=7.56"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigo_graphic_menu/js/tigo_menu_themes.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/messageclose/js/messageclose.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/detectmobilebrowser.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/jquery.wait.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/jquery.fittext.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/tigosmart_customjs.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/tigosmart_js.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_customjs/waypoints.min.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/tigosmart_custom_pages/js/panel_ajax_loader.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/field_group/field_group.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/libraries/flexslider/jquery.flexslider-min.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/flexslider/assets/js/flexslider.load.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/js/tb-megamenu-frontend.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/custom/features/display_data_set_lists_fragment/js/display_data_set_lists_fragment.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/modules/contrib/tb_megamenu/js/tb-megamenu-touch.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/themes/omega/omega/js/jquery.formalize.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/themes/omega/omega/js/omega-mediaqueries.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/themes/tigo_smart/js/jquery.mmenu.js?p5wf0x"></script>
<script type="text/javascript" src="https://www.tigo.com.sv/sites/all/themes/tigo_smart/js/tigowebcorp.scripts.js?p5wf0x"></script>
</body>
</html>