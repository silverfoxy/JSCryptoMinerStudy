<!DOCTYPE html>


<html xmlns='http://www.w3.org/1999/xhtml'>
<head>
<title>Davivienda El Salvador</title>
<meta content='ISO-8859-1' http-equiv='content-type'>
<meta content='' name='description'>
<meta content='' name='keywords'>
<link href="css/site.css" media="screen" rel="stylesheet"
	type="text/css" />
 <script type="text/javascript" src="js/DP.js" ></script>
       
    <script type="text/javascript">
		window.onload = DP.inicio;
	</script>
	<style type="text/css">
		*{padding:0;margin:0;border:0;}
	</style>








<body>
<div id='main'>
<div class='shadow-main'>
<div class='main'>
<div class='header'>
<div class='logo'><a href="/"><img
	alt="Logo-davivienda-hsbc" src="images/logo-davivienda-hsbc.png" /></a></div>
<div class='date'>
<script type="text/JavaScript" language="JavaScript">
dows = new Array("Domingo","Lunes","Martes","Mi�rcoles","Jueves","Viernes","S�bado");
months = new Array("enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre");
now = new Date();
dow = now.getDay();
d = now.getDate();
m = now.getMonth();
h = now.getTime();
y = now.getFullYear();
document.write(dows[dow] + ", " + d + " de " + months[m] + " de " + y + "");
</script>
<br>
<div align="right">
<b>
EL SALVADOR
</b>
 </div>
</div>
</div>



<!-- 
	







              <ul class='main-menu'>

                <li>
                  <a href="/?cat=8">Otros</a>
                </li>

                <li>
                  <a href="/?cat=7">Escr&iacute;banos</a>
                </li>

                <li>
                  <a href="/?cat=6">Cajeros y Agencias</a>
                </li>

                <li>
                  <a href="/?cat=5">Corporativo</a>
                </li>

                <li>
                  <a href="/?cat=4">Davivienda Empresas</a>
                </li>

                <li>
                  <a href="/?cat=3">Banca de Personas</a>
                </li>
                <li>
                  <a href="/">Inicio</a>
                </li>
              </ul>
          
 --> <!-- inicio seccion left -->
<div class='left-h'><!-- Inicio categoria -->
<h2 class='title-h'><a
	href="/?cat=3">Banca
Personas</a></h2>
<div class='item-home'>

<h3 class='stitle-h'><a
	href="/?cat=1313">Premium</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1005">Cr&eacute;ditos</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1326">Corresponsales Financieros</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1000">Tarjetas</a>
</h3>

<div class='see_servs'><a
	href="/?cat=3">m&aacute;s
servicios</a></div>
</div>


<h2 class='title-h'><a
	href="/?cat=4">Empresas</a>
</h2>
<div class='item-home'>

<h3 class='stitle-h'><a
	href="/?cat=1012">Financiamiento</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1301">Gesti&oacute;n de Cuentas</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1008">Seguros</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1011">Comercio Exterior</a>
</h3>

<div class='see_servs'><a
	href="/?cat=4">m&aacute;s
servicios</a></div>
</div>





<h2 class='title-h'><a
	href="/?cat=5">Corporativo</a>
</h2>
<div class='item-home'>

<h3 class='stitle-h'><a
	href="/?cat=1015">Financiamiento</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1018">Cuentas por Cobrar</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1019">Seguros</a>
</h3>

<h3 class='stitle-h'><a
	href="/?cat=1020">Comercio Exterior</a>
</h3>

<div class='see_servs'><a
	href="/?cat=5">m&aacute;s
servicios</a></div>
</div>



<!-- fin categoria --></div>
<!-- fin seccion left -->





<div class='center-h'>
<div class='slider-h'>
<div id='slideShow'>
<div class='item-home-pics'>
<div class='picture-home-pics'><a
	href="http://www.davivienda.com.sv/uploaded/content/category/Convenio.pdf">  <object
classid="clsid:D27CDB6E-AE6D-11cf-96B8-444553540000" 
codebase="http://download.macromedia.com
/pub/shockwave/cabs/flash/swflash.cab#version=6,0,0,0"
width="607" height="300" id="movie" align="">
<param name="movie" value="/pics/content/banner/cominicado3.swf" >
<embed src="/pics/content/banner/cominicado3.swf"  quality="high" width="607" 
height="300" name="movie" align="" 
type="application/x-shockwave-flash"
plug inspage="http://www.macromedia.com/go/getflashplayer"> 
</object>
 </a></div>
</div>
</div>
</div>
<div id='nav'></div>
<div class='clear'></div>
<div class='more-lnks'>
<div class='bannr'>

<a
	href="http://www.davivienda.com.sv/?cat=1321">
	
	<img
	alt="" src="/pics/content/banner/canalew.jpg" title="" />
	</a>
	</div>
<div class='bannr'>
<a
	href="http://www.davivienda.com.sv/?cat=1318">
	
	<img
	alt="" src="/pics/content/banner/tarjeta.jpg" title="" />
	</a>
	</div>
<div class='bannr'>
<a
	href="http://www.davivienda.com.sv/seguros">
	
	<img
	alt="" src="/pics/content/banner/seguros web.jpg" title="" />
	</a>
</div>
<div class='bannr'>
<a
	href="https://daviviendaenlinea.davivienda.com.sv:4443/CorteTarjeta/">
	
	<img
	alt="" src="/pics/content/banner/corte2.jpg" title="" />
	</a>
</div>
<div class='clear'></div>
</div>
</div>



<div class='right-h'>


<a href="/atencion"><img src="images/logo-atencion-en-linea.png" /></a>

	
	









            <div class='banca'>
              <img alt="Top-banca" class="block" src="images/top-banca.png" />
              <div class='banca-content'>
                <h2 class='title-h-no-lnk'>
                  Banca Digital
                </h2>
                <div class='banca-detail'>
                  <p>
						
								<a href="https://bancaelectronica.davivienda.com.sv/PersonalBanking/login.davivienda" target="" >Conexi&oacute;n Personal</a> <br/>
						
								<a href="https://bancaempresaplus.davivienda.com.sv" target="_blank" >Banca Empresa Plus</a> <br/>
						
								<a href="https://bancaelectronica.davivienda.com.sv/pyme" target="" >Banc@Pyme.com</a> <br/>
						
								<a href="https://empresarialmultilatina.davivienda.com" target="_blank" >Empresarial Multilatina</a> <br/>
						
								<a href="https://bancaelectronica.davivienda.com.sv/TransaccionesInterBCR/" target="_blank" >Declaraci&oacute;n de Divisas</a> <br/>
						
                  </p>
                </div>
              </div>
              <img alt="Bottom-banca" class="block" src="images/bottom-banca.png" />
            </div>
 







<h2 class='title-h'>
              <a href="#">Noticias</a>
            </h2>
            <div class='news-home'>


            
            
              <div class='see_all_link_bold'>
                <a href="/?cat=-1">Ver todas las noticias</a>
              </div>
            </div>

	
	<h2 class='title-h'>
	<a href="/?cat=1202">Activos Extraordinarios</a>
	</h2>
	

	
	<ul id="diapos">

  
   
   
       <li>
       		
      		<a href="/?cat=1202">
				<img
				src		="pics/content/inmueble/IMG_20170706_120622.jpg" width="160px" height="120px"  
				title	="Terreno de playa" 
				alt		="Terreno de playa"/>
			</a>
			<h3 class="title-picture-diapos" align="center">
				Terreno de playa
			</h3>	
		</li>
	
	


  
   
   
       <li>
       		
      		<a href="/?cat=1202">
				<img
				src		="pics/content/inmueble/Joya de las Piletas.JPG" width="160px" height="120px"  
				title	="Vivienda" 
				alt		="Vivienda"/>
			</a>
			<h3 class="title-picture-diapos" align="center">
				Vivienda
			</h3>	
		</li>
	
	


  
   
   
       <li>
       		
      		<a href="/?cat=1202">
				<img
				src		="pics/content/inmueble/Rosal.JPG" width="160px" height="120px"  
				title	="Vivienda" 
				alt		="Vivienda"/>
			</a>
			<h3 class="title-picture-diapos" align="center">
				Vivienda
			</h3>	
		</li>
	
	



</ul>

	
	
	</div>
<div class='clear'></div>
<script type="text/javascript" src="javascript/validaciones.js"></script>








          <div id='footer'>
            <div class='footer'>

              <a href="/?cat=1025">Informaci&oacute;n institucional</a>
              <span>
                |
              </span>

              <a href="/?cat=1023">Requerimientos</a>
              <span>
                |
              </span>

              <a href="/?cat=1024">Legal</a>
              <span>
                |
              </span>

              <a href="/?cat=1207">Memorias de Labores</a>
              <span>
                |
              </span>

              <a href="/?cat=1177">Modelo de Escrituraci&oacute;n</a>
              <span>
                |
              </span>

            </div>
          </div>
          
          <div id='credits'>
            <div class='credits'>
              <p>Todos los derechos reservados &reg;&nbsp; <strong>DAVIVIENDA 2014</strong></p>
            </div>
          </div>
        </div>
        <div class='shadow-bot'></div>
      </div>
    </div>
  </body>
</html>