<!DOCTYPE html>
<html lang="es-ES" prefix="og: http://ogp.me/ns#">
<head>
	<meta name="google-site-verification" content="TR-YkLp4WHYoHln9v_02kjzvZPWLnzGO-opekDS46tk" />
<meta charset="UTF-8" >
<meta name="viewport" id="viewport" content="width=device-width, initial-scale=1.0, maximum-scale=1.0, minimum-scale=1.0, user-scalable=no" />
<link rel="shortcut icon" href="/wp-content/uploads/2018/02/favicon.png" /><link rel="pingback" href="http://cronio.sv/xmlrpc.php" />
<meta property="og:description" content="El encuentro de todos los lectores de las mejores noticias." />
<title>Portada - Diario Digital Cronio de El Salvador</title>

<!-- This site is optimized with the Yoast SEO plugin v6.3.1 - https://yoast.com/wordpress/plugins/seo/ -->
<meta name="description" content="Noticias de El Salvador Diario Digital de El Salvador, Encuentra los mejores titulares nacionales y del mundo. Diario Digital Cronio es el centro de encuentro de todos los amantes a las noticias de ultima hora y en tendencia."/>
<link rel="canonical" href="http://cronio.sv/" />
<meta property="og:locale" content="es_ES" />
<meta property="og:type" content="website" />
<meta property="og:title" content="Portada - Diario Digital Cronio de El Salvador" />
<meta property="og:description" content="Noticias de El Salvador Diario Digital de El Salvador, Encuentra los mejores titulares nacionales y del mundo. Diario Digital Cronio es el centro de encuentro de todos los amantes a las noticias de ultima hora y en tendencia." />
<meta property="og:url" content="http://cronio.sv/" />
<meta property="og:site_name" content="Diario Digital Cronio de El Salvador" />
<meta name="twitter:card" content="summary_large_image" />
<meta name="twitter:description" content="Noticias de El Salvador Diario Digital de El Salvador, Encuentra los mejores titulares nacionales y del mundo. Diario Digital Cronio es el centro de encuentro de todos los amantes a las noticias de ultima hora y en tendencia." />
<meta name="twitter:title" content="Portada - Diario Digital Cronio de El Salvador" />
<script type='application/ld+json'>{"@context":"http:\/\/schema.org","@type":"WebSite","@id":"#website","url":"http:\/\/cronio.sv\/","name":"Diario Digital Cronio de El Salvador","potentialAction":{"@type":"SearchAction","target":"http:\/\/cronio.sv\/?s={search_term_string}","query-input":"required name=search_term_string"}}</script>
<!-- / Yoast SEO plugin. -->

<link rel='dns-prefetch' href='//fonts.googleapis.com' />
<link rel='dns-prefetch' href='//s.w.org' />
<link rel="alternate" type="application/rss+xml" title="Diario Digital Cronio de El Salvador &raquo; Feed" href="http://cronio.sv/feed/" />
<link rel="alternate" type="application/rss+xml" title="Diario Digital Cronio de El Salvador &raquo; RSS de los comentarios" href="http://cronio.sv/comments/feed/" />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/cronio.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.9.4"}};
			!function(a,b,c){function d(a,b){var c=String.fromCharCode;l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,a),0,0);var d=k.toDataURL();l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,b),0,0);var e=k.toDataURL();return d===e}function e(a){var b;if(!l||!l.fillText)return!1;switch(l.textBaseline="top",l.font="600 32px Arial",a){case"flag":return!(b=d([55356,56826,55356,56819],[55356,56826,8203,55356,56819]))&&(b=d([55356,57332,56128,56423,56128,56418,56128,56421,56128,56430,56128,56423,56128,56447],[55356,57332,8203,56128,56423,8203,56128,56418,8203,56128,56421,8203,56128,56430,8203,56128,56423,8203,56128,56447]),!b);case"emoji":return b=d([55357,56692,8205,9792,65039],[55357,56692,8203,9792,65039]),!b}return!1}function f(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var g,h,i,j,k=b.createElement("canvas"),l=k.getContext&&k.getContext("2d");for(j=Array("flag","emoji"),c.supports={everything:!0,everythingExceptFlag:!0},i=0;i<j.length;i++)c.supports[j[i]]=e(j[i]),c.supports.everything=c.supports.everything&&c.supports[j[i]],"flag"!==j[i]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[j[i]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(h=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",h,!1),a.addEventListener("load",h,!1)):(a.attachEvent("onload",h),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),g=c.source||{},g.concatemoji?f(g.concatemoji):g.wpemoji&&g.twemoji&&(f(g.twemoji),f(g.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='stylesheet' id='svc-font-awesome-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-team/../assets/css/font-awesome.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='svc-hover-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-team/../assets/css/hover.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='mvp-custom-style-css'  href='http://cronio.sv/wp-content/themes/zox-news/style.css?ver=4.9.4' type='text/css' media='all' />
<style id='mvp-custom-style-inline-css' type='text/css'>


#mvp-wallpaper {
	background: url() no-repeat 50% 0;
	}

#mvp-foot-copy a {
	color: #0be6af;
	}

#mvp-content-main p a,
.mvp-post-add-main p a {
	box-shadow: inset 0 -4px 0 #0be6af;
	}

#mvp-content-main p a:hover,
.mvp-post-add-main p a:hover {
	background: #0be6af;
	}

a,
a:visited,
.post-info-name a,
.woocommerce .woocommerce-breadcrumb a {
	color: #c93639;
	}

#mvp-side-wrap a:hover {
	color: #c93639;
	}

.mvp-fly-top:hover,
.mvp-vid-box-wrap,
ul.mvp-soc-mob-list li.mvp-soc-mob-com {
	background: #c93639;
	}

nav.mvp-fly-nav-menu ul li.menu-item-has-children:after,
.mvp-feat1-left-wrap span.mvp-cd-cat,
.mvp-widget-feat1-top-story span.mvp-cd-cat,
.mvp-widget-feat2-left-cont span.mvp-cd-cat,
.mvp-widget-dark-feat span.mvp-cd-cat,
.mvp-widget-dark-sub span.mvp-cd-cat,
.mvp-vid-wide-text span.mvp-cd-cat,
.mvp-feat2-top-text span.mvp-cd-cat,
.mvp-feat3-main-story span.mvp-cd-cat,
.mvp-feat3-sub-text span.mvp-cd-cat,
.mvp-feat4-main-text span.mvp-cd-cat,
.woocommerce-message:before,
.woocommerce-info:before,
.woocommerce-message:before {
	color: #c93639;
	}

#searchform input,
.mvp-authors-name {
	border-bottom: 1px solid #c93639;
	}

.mvp-fly-top:hover {
	border-top: 1px solid #c93639;
	border-left: 1px solid #c93639;
	border-bottom: 1px solid #c93639;
	}

.woocommerce .widget_price_filter .ui-slider .ui-slider-handle,
.woocommerce #respond input#submit.alt,
.woocommerce a.button.alt,
.woocommerce button.button.alt,
.woocommerce input.button.alt,
.woocommerce #respond input#submit.alt:hover,
.woocommerce a.button.alt:hover,
.woocommerce button.button.alt:hover,
.woocommerce input.button.alt:hover {
	background-color: #c93639;
	}

.woocommerce-error,
.woocommerce-info,
.woocommerce-message {
	border-top-color: #c93639;
	}

ul.mvp-feat1-list-buts li.active span.mvp-feat1-list-but,
span.mvp-widget-home-title,
span.mvp-post-cat,
span.mvp-feat1-pop-head {
	background: #c93639;
	}

.woocommerce span.onsale {
	background-color: #c93639;
	}

.mvp-widget-feat2-side-more-but,
.woocommerce .star-rating span:before,
span.mvp-prev-next-label,
.mvp-cat-date-wrap .sticky {
	color: #c93639 !important;
	}

#mvp-main-nav-top,
#mvp-fly-wrap,
.mvp-soc-mob-right,
#mvp-main-nav-small-cont {
	background: #000000;
	}

#mvp-main-nav-small .mvp-fly-but-wrap span,
#mvp-main-nav-small .mvp-search-but-wrap span,
.mvp-nav-top-left .mvp-fly-but-wrap span,
#mvp-fly-wrap .mvp-fly-but-wrap span {
	background: #555555;
	}

.mvp-nav-top-right .mvp-nav-search-but,
span.mvp-fly-soc-head,
.mvp-soc-mob-right i,
#mvp-main-nav-small span.mvp-nav-search-but,
#mvp-main-nav-small .mvp-nav-menu ul li a  {
	color: #555555;
	}

#mvp-main-nav-small .mvp-nav-menu ul li.menu-item-has-children a:after {
	border-color: #555555 transparent transparent transparent;
	}

#mvp-nav-top-wrap span.mvp-nav-search-but:hover,
#mvp-main-nav-small span.mvp-nav-search-but:hover {
	color: #0be6af;
	}

#mvp-nav-top-wrap .mvp-fly-but-wrap:hover span,
#mvp-main-nav-small .mvp-fly-but-wrap:hover span,
span.mvp-woo-cart-num:hover {
	background: #0be6af;
	}

#mvp-main-nav-bot-cont {
	background: #ffffff;
	}

#mvp-nav-bot-wrap .mvp-fly-but-wrap span,
#mvp-nav-bot-wrap .mvp-search-but-wrap span {
	background: #000000;
	}

#mvp-nav-bot-wrap span.mvp-nav-search-but,
#mvp-nav-bot-wrap .mvp-nav-menu ul li a {
	color: #000000;
	}

#mvp-nav-bot-wrap .mvp-nav-menu ul li.menu-item-has-children a:after {
	border-color: #000000 transparent transparent transparent;
	}

.mvp-nav-menu ul li:hover a {
	border-bottom: 5px solid #c93639;
	}

#mvp-nav-bot-wrap .mvp-fly-but-wrap:hover span {
	background: #c93639;
	}

#mvp-nav-bot-wrap span.mvp-nav-search-but:hover {
	color: #c93639;
	}

body,
.mvp-feat1-feat-text p,
.mvp-feat2-top-text p,
.mvp-feat3-main-text p,
.mvp-feat3-sub-text p,
#searchform input,
.mvp-author-info-text,
span.mvp-post-excerpt,
.mvp-nav-menu ul li ul.sub-menu li a,
nav.mvp-fly-nav-menu ul li a,
.mvp-ad-label,
span.mvp-feat-caption,
.mvp-post-tags a,
.mvp-post-tags a:visited,
span.mvp-author-box-name a,
#mvp-author-box-text p,
.mvp-post-gallery-text p,
ul.mvp-soc-mob-list li span,
#comments,
h3#reply-title,
h2.comments,
#mvp-foot-copy p,
span.mvp-fly-soc-head,
.mvp-post-tags-header,
span.mvp-prev-next-label,
span.mvp-post-add-link-but,
#mvp-comments-button a,
#mvp-comments-button span.mvp-comment-but-text,
.woocommerce ul.product_list_widget span.product-title,
.woocommerce ul.product_list_widget li a,
.woocommerce #reviews #comments ol.commentlist li .comment-text p.meta,
.woocommerce div.product p.price,
.woocommerce div.product p.price ins,
.woocommerce div.product p.price del,
.woocommerce ul.products li.product .price del,
.woocommerce ul.products li.product .price ins,
.woocommerce ul.products li.product .price,
.woocommerce #respond input#submit,
.woocommerce a.button,
.woocommerce button.button,
.woocommerce input.button,
.woocommerce .widget_price_filter .price_slider_amount .button,
.woocommerce span.onsale,
.woocommerce-review-link,
#woo-content p.woocommerce-result-count,
.woocommerce div.product .woocommerce-tabs ul.tabs li a,
a.mvp-inf-more-but,
span.mvp-cont-read-but,
span.mvp-cd-cat,
span.mvp-cd-date,
.mvp-feat4-main-text p,
span.mvp-woo-cart-num,
span.mvp-widget-home-title2,
.wp-caption,
#mvp-content-main p.wp-caption-text,
.gallery-caption,
.mvp-post-add-main p.wp-caption-text,
#bbpress-forums,
#bbpress-forums p,
.protected-post-form input,
#mvp-feat6-text p {
	font-family: 'Arial', sans-serif;
	}

.mvp-blog-story-text p,
span.mvp-author-page-desc,
#mvp-404 p,
.mvp-widget-feat1-bot-text p,
.mvp-widget-feat2-left-text p,
.mvp-flex-story-text p,
.mvp-search-text p,
#mvp-content-main p,
.mvp-post-add-main p,
.rwp-summary,
.rwp-u-review__comment,
.mvp-feat5-mid-main-text p,
.mvp-feat5-small-main-text p {
	font-family: 'PT Serif', sans-serif;
	}

.mvp-nav-menu ul li a,
#mvp-foot-menu ul li a {
	font-family: 'Oswald', sans-serif;
	}


.mvp-feat1-sub-text h2,
.mvp-feat1-pop-text h2,
.mvp-feat1-list-text h2,
.mvp-widget-feat1-top-text h2,
.mvp-widget-feat1-bot-text h2,
.mvp-widget-dark-feat-text h2,
.mvp-widget-dark-sub-text h2,
.mvp-widget-feat2-left-text h2,
.mvp-widget-feat2-right-text h2,
.mvp-blog-story-text h2,
.mvp-flex-story-text h2,
.mvp-vid-wide-more-text p,
.mvp-prev-next-text p,
.mvp-related-text,
.mvp-post-more-text p,
h2.mvp-authors-latest a,
.mvp-feat2-bot-text h2,
.mvp-feat3-sub-text h2,
.mvp-feat3-main-text h2,
.mvp-feat4-main-text h2,
.mvp-feat5-text h2,
.mvp-feat5-mid-main-text h2,
.mvp-feat5-small-main-text h2,
.mvp-feat5-mid-sub-text h2,
#mvp-feat6-text h2 {
	font-family: 'Oswald', sans-serif;
	}

.mvp-feat2-top-text h2,
.mvp-feat1-feat-text h2,
h1.mvp-post-title,
h1.mvp-post-title-wide,
.mvp-drop-nav-title h4,
#mvp-content-main blockquote p,
.mvp-post-add-main blockquote p,
#mvp-404 h1,
#woo-content h1.page-title,
.woocommerce div.product .product_title,
.woocommerce ul.products li.product h3 {
	font-family: 'Arial', sans-serif;
	}

span.mvp-feat1-pop-head,
.mvp-feat1-pop-text:before,
span.mvp-feat1-list-but,
span.mvp-widget-home-title,
.mvp-widget-feat2-side-more,
span.mvp-post-cat,
span.mvp-page-head,
h1.mvp-author-top-head,
.mvp-authors-name,
#mvp-content-main h1,
#mvp-content-main h2,
#mvp-content-main h3,
#mvp-content-main h4,
#mvp-content-main h5,
#mvp-content-main h6,
.woocommerce .related h2,
.woocommerce div.product .woocommerce-tabs .panel h2,
.woocommerce div.product .product_title,
.mvp-feat5-side-list .mvp-feat1-list-img:after {
	font-family: 'Arial', sans-serif;
	}

	

	.mvp-vid-box-wrap,
	.mvp-feat1-left-wrap span.mvp-cd-cat,
	.mvp-widget-feat1-top-story span.mvp-cd-cat,
	.mvp-widget-feat2-left-cont span.mvp-cd-cat,
	.mvp-widget-dark-feat span.mvp-cd-cat,
	.mvp-widget-dark-sub span.mvp-cd-cat,
	.mvp-vid-wide-text span.mvp-cd-cat,
	.mvp-feat2-top-text span.mvp-cd-cat,
	.mvp-feat3-main-story span.mvp-cd-cat {
		color: #fff;
		}
		

	#mvp-main-nav-top {
		background: #fff;
		padding: 15px 0 0;
		}
	#mvp-fly-wrap,
	.mvp-soc-mob-right,
	#mvp-main-nav-small-cont {
		background: #fff;
		}
	#mvp-main-nav-small .mvp-fly-but-wrap span,
	#mvp-main-nav-small .mvp-search-but-wrap span,
	.mvp-nav-top-left .mvp-fly-but-wrap span,
	#mvp-fly-wrap .mvp-fly-but-wrap span {
		background: #000;
		}
	.mvp-nav-top-right .mvp-nav-search-but,
	span.mvp-fly-soc-head,
	.mvp-soc-mob-right i,
	#mvp-main-nav-small span.mvp-nav-search-but,
	#mvp-main-nav-small .mvp-nav-menu ul li a  {
		color: #000;
		}
	#mvp-main-nav-small .mvp-nav-menu ul li.menu-item-has-children a:after {
		border-color: #000 transparent transparent transparent;
		}
	.mvp-feat1-feat-text h2,
	h1.mvp-post-title,
	.mvp-feat2-top-text h2,
	.mvp-feat3-main-text h2,
	#mvp-content-main blockquote p,
	.mvp-post-add-main blockquote p {
		font-family: 'Anton', sans-serif;
		font-weight: 400;
		letter-spacing: normal;
		}
	.mvp-feat1-feat-text h2,
	.mvp-feat2-top-text h2,
	.mvp-feat3-main-text h2 {
		line-height: 1;
		text-transform: uppercase;
		}
		

	span.mvp-nav-soc-but,
	ul.mvp-fly-soc-list li a,
	span.mvp-woo-cart-num {
		background: rgba(0,0,0,.8);
		}
	span.mvp-woo-cart-icon {
		color: rgba(0,0,0,.8);
		}
	nav.mvp-fly-nav-menu ul li,
	nav.mvp-fly-nav-menu ul li ul.sub-menu {
		border-top: 1px solid rgba(0,0,0,.1);
		}
	nav.mvp-fly-nav-menu ul li a {
		color: #000;
		}
	.mvp-drop-nav-title h4 {
		color: #000;
		}
		

	.mvp-nav-links {
		display: none;
		}
		
</style>
<link rel='stylesheet' id='mvp-reset-css'  href='http://cronio.sv/wp-content/themes/zox-news/css/reset.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='fontawesome-css'  href='http://cronio.sv/wp-content/themes/zox-news/font-awesome/css/font-awesome.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='mvp-fonts-css'  href='//fonts.googleapis.com/css?family=Advent+Pro%3A700%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7COpen+Sans%3A700%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7CAnton%3A400%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7COswald%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7CArial%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7CArial%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7CArial%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7CPT+Serif%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese%7COswald%3A100%2C200%2C300%2C400%2C500%2C600%2C700%2C800%2C900%26subset%3Dlatin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek-ext%2Cgreek%2Cvietnamese' type='text/css' media='all' />
<link rel='stylesheet' id='mvp-media-queries-css'  href='http://cronio.sv/wp-content/themes/zox-news/css/media-queries.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='svc-imagehover-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc/../assets/css/imagehover.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='svc-justifiedGallery-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc/../assets/css/justifiedGallery.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='svc-megnific-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/css/magnific-popup.css?ver=4.9.4' type='text/css' media='all' />
<script type='text/javascript' src='http://cronio.sv/wp-includes/js/jquery/jquery.js?ver=1.12.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-includes/js/jquery/jquery-migrate.min.js?ver=1.4.1'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/js/isotope.pkgd.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-soc/../assets/js/jquery.viewportchecker.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-soc/../assets/js/doT.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-soc/../assets/js/moment-with-locales.min.js?ver=4.9.4'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var svc_ajax_url = {"url":"http:\/\/cronio.sv\/wp-admin\/admin-ajax.php","laungage":"es_ES"};
/* ]]> */
</script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-soc/../assets/js/social-stream.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/js/megnific.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc/../assets/js/jquery.justifiedGallery.min.js?ver=4.9.4'></script>
<link rel='https://api.w.org/' href='http://cronio.sv/wp-json/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://cronio.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://cronio.sv/wp-includes/wlwmanifest.xml" /> 
<link rel='shortlink' href='http://cronio.sv/' />
<link rel="alternate" type="application/json+oembed" href="http://cronio.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fcronio.sv%2F" />
<link rel="alternate" type="text/xml+oembed" href="http://cronio.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fcronio.sv%2F&#038;format=xml" />

<!-- This site is using AdRotate v4.9 to display their advertisements - https://ajdg.solutions/products/adrotate-for-wordpress/ -->
<!-- AdRotate CSS -->
<style type="text/css" media="screen">
	.g { margin:0px; padding:0px; overflow:hidden; line-height:1; zoom:1; }
	.g img { height:auto; }
	.g-col { position:relative; float:left; }
	.g-col:first-child { margin-left: 0; }
	.g-col:last-child { margin-right: 0; }
	.g-1 { margin:0px;width:100%; max-width:300px; height:100%; max-height:250px; }
	@media only screen and (max-width: 480px) {
		.g-col, .g-dyn, .g-single { width:100%; margin-left:0; margin-right:0; }
	}
</style>
<!-- /AdRotate CSS -->

    <style>
	.svc_post_grid_list_container{ display:none;}
	#loader {background-image: url("http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc/../assets/css/loader.GIF");}
	</style>
        <style>
	.svc_social_stream_container{ display:none;}
	#loader {background-image: url("http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-soc/../assets/css/loader.GIF");}
	</style>
        <style>
	.svc_post_grid_list_container{ display:none;}
	#loader {background-image: url("http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/css/loader.GIF");}
	</style>
        <style>
	.svc_post_grid_list_container{ display:none;}
	#loader {background-image: url("http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-post/../assets/css/loader.GIF");}
	</style>
    		<style type="text/css">.recentcomments a{display:inline !important;padding:0 !important;margin:0 !important;}</style>
		</head>
<body class="home page-template page-template-page-home page-template-page-home-php page page-id-17">
	<!-- Start Alexa AMP Certify Javascript -->
<amp-analytics type="alexametrics">
<script type="application/json"> {"vars": { "atrk_acct": "2bRCo1IWhe105T", "domain": "cronio.sv" }}</script>
</amp-analytics>
<!-- End Alexa AMP Certify Javascript -->   
	<div id="mvp-fly-wrap">
	<div id="mvp-fly-menu-top" class="left relative">
		<div class="mvp-fly-top-out left relative">
			<div class="mvp-fly-top-in">
				<div id="mvp-fly-logo" class="left relative">
											<a href="http://cronio.sv/"><img src="http://cronio.sv/wp-content/uploads/2018/03/BANNERHOMECRONIO-1.png" alt="Diario Digital Cronio de El Salvador" data-rjs="2" /></a>
									</div><!--mvp-fly-logo-->
			</div><!--mvp-fly-top-in-->
			<div class="mvp-fly-but-wrap mvp-fly-but-menu mvp-fly-but-click">
				<span></span>
				<span></span>
				<span></span>
				<span></span>
			</div><!--mvp-fly-but-wrap-->
		</div><!--mvp-fly-top-out-->
	</div><!--mvp-fly-menu-top-->
	<div id="mvp-fly-menu-wrap">
		<nav class="mvp-fly-nav-menu left relative">
			<div class="menu-principal-container"><ul id="menu-principal" class="menu"><li id="menu-item-20" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-home current-menu-item page_item page-item-17 current_page_item menu-item-20"><a href="http://cronio.sv/">Portada</a></li>
<li id="menu-item-8" class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-8"><a href="http://cronio.sv/category/nacionales/">Nacionales</a></li>
<li id="menu-item-14" class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-14"><a href="http://cronio.sv/category/politica/">Política</a></li>
<li id="menu-item-9" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-9"><a href="http://cronio.sv/category/internacionales/">Internacionales</a></li>
<li id="menu-item-12" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-12"><a href="http://cronio.sv/category/negocios/">Negocios</a></li>
<li id="menu-item-11" class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-11"><a href="http://cronio.sv/category/deportes/">Deportes</a></li>
<li id="menu-item-10" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-10"><a href="http://cronio.sv/category/croniotv/">CronioTV</a></li>
<li id="menu-item-16" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-16"><a href="http://cronio.sv/category/tendencias/">Tendencias</a></li>
<li id="menu-item-13" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-13"><a href="http://cronio.sv/category/opinet/">Opinet</a></li>
<li id="menu-item-15" class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-15"><a href="http://cronio.sv/category/redes/">Redes</a></li>
</ul></div>		</nav>
	</div><!--mvp-fly-menu-wrap-->
	<div id="mvp-fly-soc-wrap">
		<span class="mvp-fly-soc-head">Connect with us</span>
		<ul class="mvp-fly-soc-list left relative">
							<li><a href="https://www.facebook.com/croniosv/" target="_blank" class="fa fa-facebook fa-2"></a></li>
										<li><a href="https://twitter.com/croniosv" target="_blank" class="fa fa-twitter fa-2"></a></li>
													<li><a href="https://www.instagram.com/croniosv/" target="_blank" class="fa fa-instagram fa-2"></a></li>
													<li><a href="https://www.youtube.com/channel/UC9uaphREcIxCZHQgmoxkn0g/videos?disable_polymer=1" target="_blank" class="fa fa-youtube-play fa-2"></a></li>
											</ul>
	</div><!--mvp-fly-soc-wrap-->
</div><!--mvp-fly-wrap-->	<div id="mvp-site" class="left relative">
		<div id="mvp-search-wrap">
			<div id="mvp-search-box">
				<form method="get" id="searchform" action="http://cronio.sv/">
	<input type="text" name="s" id="s" value="Search" onfocus='if (this.value == "Search") { this.value = ""; }' onblur='if (this.value == "") { this.value = "Search"; }' />
	<input type="hidden" id="searchsubmit" value="Search" />
</form>			</div><!--mvp-search-box-->
			<div class="mvp-search-but-wrap mvp-search-click">
				<span></span>
				<span></span>
			</div><!--mvp-search-but-wrap-->
		</div><!--mvp-search-wrap-->
				<div id="mvp-site-wall" class="left relative">
											<div id="mvp-leader-wrap">
					<a href="http://www.megablock.com.sv/"><img src="/wp-content/uploads/2018/02/megablock.jpeg" ></a>				</div><!--mvp-leader-wrap-->
										<div id="mvp-site-main" class="left relative">
			<header id="mvp-main-head-wrap" class="left relative">
									<nav id="mvp-main-nav-wrap" class="left relative">
						<div id="mvp-main-nav-top" class="left relative">
							<div class="mvp-main-box">
								<div id="mvp-nav-top-wrap" class="left relative">
									<div class="mvp-nav-top-right-out left relative">
										<div class="mvp-nav-top-right-in">
											<div class="mvp-nav-top-cont left relative">
												<div class="mvp-nav-top-left-out relative">
													<div class="mvp-nav-top-left">
														<div class="mvp-nav-soc-wrap">
																															<a href="https://www.facebook.com/croniosv/" target="_blank"><span class="mvp-nav-soc-but fa fa-facebook fa-2"></span></a>
																																														<a href="https://twitter.com/croniosv" target="_blank"><span class="mvp-nav-soc-but fa fa-twitter fa-2"></span></a>
																																														<a href="https://www.instagram.com/croniosv/" target="_blank"><span class="mvp-nav-soc-but fa fa-instagram fa-2"></span></a>
																																														<a href="https://www.youtube.com/channel/UC9uaphREcIxCZHQgmoxkn0g/videos?disable_polymer=1" target="_blank"><span class="mvp-nav-soc-but fa fa-youtube-play fa-2"></span></a>
																													</div><!--mvp-nav-soc-wrap-->
														<div class="mvp-fly-but-wrap mvp-fly-but-click left relative">
															<span></span>
															<span></span>
															<span></span>
															<span></span>
														</div><!--mvp-fly-but-wrap-->
													</div><!--mvp-nav-top-left-->
													<div class="mvp-nav-top-left-in">
														<div class="mvp-nav-top-mid left relative" itemscope itemtype="http://schema.org/Organization">
																															<a class="mvp-nav-logo-reg" itemprop="url" href="http://cronio.sv/"><img itemprop="logo" src="http://cronio.sv/wp-content/uploads/2018/03/BANNERHOMECRONIO.png" alt="Diario Digital Cronio de El Salvador" data-rjs="2" /></a>
																																														<a class="mvp-nav-logo-small" href="http://cronio.sv/"><img src="http://cronio.sv/wp-content/uploads/2018/03/BANNERHOMECRONIO-1.png" alt="Diario Digital Cronio de El Salvador" data-rjs="2" /></a>
																																														<h1 class="mvp-logo-title">Diario Digital Cronio de El Salvador</h1>
																																												</div><!--mvp-nav-top-mid-->
													</div><!--mvp-nav-top-left-in-->
												</div><!--mvp-nav-top-left-out-->
											</div><!--mvp-nav-top-cont-->
										</div><!--mvp-nav-top-right-in-->
										<div class="mvp-nav-top-right">
																						<span class="mvp-nav-search-but fa fa-search fa-2 mvp-search-click"></span>
										</div><!--mvp-nav-top-right-->
									</div><!--mvp-nav-top-right-out-->
								</div><!--mvp-nav-top-wrap-->
							</div><!--mvp-main-box-->
						</div><!--mvp-main-nav-top-->
						<div id="mvp-main-nav-bot" class="left relative">
							<div id="mvp-main-nav-bot-cont" class="left">
								<div class="mvp-main-box">
									<div id="mvp-nav-bot-wrap" class="left">
										<div class="mvp-nav-bot-right-out left">
											<div class="mvp-nav-bot-right-in">
												<div class="mvp-nav-bot-cont left">
													<div class="mvp-nav-bot-left-out">
														<div class="mvp-nav-bot-left left relative">
															<div class="mvp-fly-but-wrap mvp-fly-but-click left relative">
																<span></span>
																<span></span>
																<span></span>
																<span></span>
															</div><!--mvp-fly-but-wrap-->
														</div><!--mvp-nav-bot-left-->
														<div class="mvp-nav-bot-left-in">
															<div class="mvp-nav-menu left">
																<div class="menu-principal-container"><ul id="menu-principal-1" class="menu"><li class="menu-item menu-item-type-post_type menu-item-object-page menu-item-home current-menu-item page_item page-item-17 current_page_item menu-item-20"><a href="http://cronio.sv/">Portada</a></li>
<li class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-8"><a href="http://cronio.sv/category/nacionales/">Nacionales</a><div class="mvp-mega-dropdown"><div class="mvp-main-box"><ul class="mvp-mega-list"><li><a href="http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/esposados-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/esposados-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/esposados-300x180.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/esposados-768x462.jpg 768w, http://cronio.sv/wp-content/uploads/2018/03/esposados-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/esposados.jpg 900w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Investigadores de la PNC son capturados por matar a otro agente y alterar la escena del crimen</p></a></li><li><a href="http://cronio.sv/nacionales/pnc-captura-14-pandilleros-ahuachapan/"><div class="mvp-mega-img"><img width="400" height="211" src="http://cronio.sv/wp-content/uploads/2018/03/DYw8zE_WAAAzl2R-400x211.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" /></div><p>PNC captura a 14 pandilleros en Ahuachapán </p></a></li><li><a href="http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Juez ordena que Jorge Hernández, conciliara con algunos periodistas a quienes habría retenido cuotas de Seguro Social y AFP</p></a></li><li><a href="http://cronio.sv/nacionales/bulevar-venezuela-cerrado-accidente-transito/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521586878-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521586878-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521586878-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Bulevar Venezuela cerrado por accidente de tránsito</p></a></li><li><a href="http://cronio.sv/nacionales/pnc-captura-medico-quien-acusado-abusar-una-joven-usulutan/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521575580-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521575580-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521575580-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>PNC captura a Medico quien es acusado de abusar de una joven en Usulután</p></a></li></ul></div></div></li>
<li class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-14"><a href="http://cronio.sv/category/politica/">Política</a><div class="mvp-mega-dropdown"><div class="mvp-main-box"><ul class="mvp-mega-list"><li><a href="http://cronio.sv/politica/carlos-caceres-anuncia-sera-nuevo-embajador-mexico/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Carlos Cáceres, anuncia que sera el nuevo Embajador en México</p></a></li><li><a href="http://cronio.sv/politica/lopez-davidson-cambios-gobierno-fue-reciclaje-decorativo-los-mismos-funcionarios/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tavo-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tavo-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/tavo-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>López Davidson: &#8220;Cambios en el Gobierno fue un reciclaje decorativo de los mismos funcionarios&#8221;</p></a></li><li><a href="http://cronio.sv/politica/smartmatic-sera-demanda-tse-confirma-julio-olivo/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Smartmatic será demanda por el TSE confirma Julio Olivo</p></a></li><li><a href="http://cronio.sv/politica/ya-no-habran-mas-cambios-gabinete-gobierno-dice-roberto-lorenzana/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Ya no habrán más cambios en el gabinete de gobierno dice Roberto Lorenzana</p></a></li><li><a href="http://cronio.sv/politica/norman-quijano-aspira-la-presidencia-la-asamblea-legislativa-gracias-al-voto-popular/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Norman Quijano aspira a la presidencia de la Asamblea Legislativa gracias al voto popular</p></a></li></ul></div></div></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-9"><a href="http://cronio.sv/category/internacionales/">Internacionales</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-12"><a href="http://cronio.sv/category/negocios/">Negocios</a></li>
<li class="mvp-mega-dropdown menu-item menu-item-type-taxonomy menu-item-object-category menu-item-11"><a href="http://cronio.sv/category/deportes/">Deportes</a><div class="mvp-mega-dropdown"><div class="mvp-main-box"><ul class="mvp-mega-list"><li><a href="http://cronio.sv/deportes/internacionales-deportes/messi-luce-la-nueva-indumentaria-alternativa-argentina-mundial-rusia-2018/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Messi luce la nueva indumentaria alternativa de Argentina para el Mundial Rusia 2018</p></a></li><li><a href="http://cronio.sv/deportes/internacionales-deportes/cristiano-ronaldo-no-nadie-mejor/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>Cristiano Ronaldo: “No hay nadie mejor que yo”</p></a></li><li><a href="http://cronio.sv/deportes/real-madrid-arrolla-al-girona-6-3/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/madrid-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/madrid-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/madrid-300x180.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/madrid-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/madrid.jpg 700w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>El Real Madrid arrolla al Girona 6-3</p></a></li><li><a href="http://cronio.sv/deportes/barca-se-impone-2-0-al-athletic-avanza-la-liga/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/barca-1-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/barca-1-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/barca-1-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>El Barca se impone 2-0 al Athletic y avanza en la Liga</p></a></li><li><a href="http://cronio.sv/deportes/messi-baila-celebrar-gol-frente-al-athletic/"><div class="mvp-mega-img"><img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/messi-400x240.jpg" class="attachment-mvp-mid-thumb size-mvp-mid-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/messi-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/messi-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/messi-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" /></div><p>VIDEO Messi baila para celebrar su gol frente al Athletic</p></a></li></ul></div></div></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-10"><a href="http://cronio.sv/category/croniotv/">CronioTV</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-16"><a href="http://cronio.sv/category/tendencias/">Tendencias</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-13"><a href="http://cronio.sv/category/opinet/">Opinet</a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-15"><a href="http://cronio.sv/category/redes/">Redes</a></li>
</ul></div>															</div><!--mvp-nav-menu-->
														</div><!--mvp-nav-bot-left-in-->
													</div><!--mvp-nav-bot-left-out-->
												</div><!--mvp-nav-bot-cont-->
											</div><!--mvp-nav-bot-right-in-->
											<div class="mvp-nav-bot-right left relative">
												<span class="mvp-nav-search-but fa fa-search fa-2 mvp-search-click"></span>
											</div><!--mvp-nav-bot-right-->
										</div><!--mvp-nav-bot-right-out-->
									</div><!--mvp-nav-bot-wrap-->
								</div><!--mvp-main-nav-bot-cont-->
							</div><!--mvp-main-box-->
						</div><!--mvp-main-nav-bot-->
					</nav><!--mvp-main-nav-wrap-->
							</header><!--mvp-main-head-wrap-->
			<div id="mvp-main-body-wrap" class="left relative">	<div class="svc_post_grid_block ">
		<div class="svc_mask " id="svc_mask_740">
			<div id="loader"></div>
		</div>

		<div class="sa_block_wrap sa_block_big_grid_1 sa-grid-style-1 sa-hover-1 " id="svc_post_grid_list_container_740">
		<div class="sa_block_inner">
			<div class="sa-big-grid-post-0 sa-big-grid-post sa-big-thumb">
				<div class="svc_share">                            
		<i class="fa fa-share-alt"></i>
		<div class="svc_share-box full-color">
		  <ul class="s8-social">
			<li class="facebook">
				<a href="https://www.facebook.com/sharer/sharer.php?u=http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/" target="_blank" title="">
					<i class="fa fa-facebook"></i>
				</a>
			</li>
			<li class="google">
				<a href="https://plusone.google.com/share?url=http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/" target="_blank" title="">
					<i class="fa fa-google-plus"></i>
				</a>
			</li>
			<li class="twitter">
				<a href="https://twitter.com/intent/tweet?text=&amp;url=http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/" target="_blank" title="">
					<i class="fa fa-twitter"></i>
				</a>
			</li>
		  </ul>
		</div>
	</div>
				<div class="sa-module-thumb">
				<a href="http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/" target="_self">
					<img width="900" height="541" src="http://cronio.sv/wp-content/uploads/2018/03/esposados.jpg" class="entry-thumb" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/esposados.jpg 900w, http://cronio.sv/wp-content/uploads/2018/03/esposados-300x180.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/esposados-768x462.jpg 768w, http://cronio.sv/wp-content/uploads/2018/03/esposados-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/esposados-400x240.jpg 400w" sizes="(max-width: 900px) 100vw, 900px" />				</a>
			</div>
			<div class="sa-meta-info-container">
				<div class="sa-meta-align">
					<div class="sa-big-grid-meta">
					<div class="svc_port_cat"><a>Judicial</a></div>						
						<h3 class="entry-title sa-module-title">
							<a href="http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/">Investigadores de la PNC son capturados por matar a otro agente y alterar la escena del crimen</a>
						</h3>
					</div>
				</div>
			</div>
		</div>
				
				
				<div class="sa-big-grid-scroll">
				<div class="sa-big-grid-post-1 sa-big-grid-post sa-small-thumb">
						<div class="svc_share">                            
		<i class="fa fa-share-alt"></i>
		<div class="svc_share-box full-color">
		  <ul class="s8-social">
			<li class="facebook">
				<a href="https://www.facebook.com/sharer/sharer.php?u=http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/" target="_blank" title="">
					<i class="fa fa-facebook"></i>
				</a>
			</li>
			<li class="google">
				<a href="https://plusone.google.com/share?url=http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/" target="_blank" title="">
					<i class="fa fa-google-plus"></i>
				</a>
			</li>
			<li class="twitter">
				<a href="https://twitter.com/intent/tweet?text=&amp;url=http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/" target="_blank" title="">
					<i class="fa fa-twitter"></i>
				</a>
			</li>
		  </ul>
		</div>
	</div>
						<div class="sa-module-thumb">
						<a href="http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/" target="_self">
							<img width="900" height="506" src="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7.jpg" class="entry-thumb" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7.jpg 900w, http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-300x169.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-768x432.jpg 768w" sizes="(max-width: 900px) 100vw, 900px" />						</a>
					</div>
					<div class="sa-meta-info-container">
						<div class="sa-meta-align">
							<div class="sa-big-grid-meta">
								<div class="svc_port_cat"><a>Judicial</a></div>								<h3 class="entry-title sa-module-title"><a href="http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/">Juez ordena que Jorge Hernández, conciliara con algunos periodistas a quienes habría retenido cuotas de Seguro Social y AFP</a></h3>
							</div>
						</div>
					</div>
				</div>
					
						<div class="sa-big-grid-post-1 sa-big-grid-post sa-small-thumb">
						<div class="svc_share">                            
		<i class="fa fa-share-alt"></i>
		<div class="svc_share-box full-color">
		  <ul class="s8-social">
			<li class="facebook">
				<a href="https://www.facebook.com/sharer/sharer.php?u=http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/" target="_blank" title="">
					<i class="fa fa-facebook"></i>
				</a>
			</li>
			<li class="google">
				<a href="https://plusone.google.com/share?url=http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/" target="_blank" title="">
					<i class="fa fa-google-plus"></i>
				</a>
			</li>
			<li class="twitter">
				<a href="https://twitter.com/intent/tweet?text=&amp;url=http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/" target="_blank" title="">
					<i class="fa fa-twitter"></i>
				</a>
			</li>
		  </ul>
		</div>
	</div>
						<div class="sa-module-thumb">
						<a href="http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/" target="_self">
							<img width="942" height="402" src="http://cronio.sv/wp-content/uploads/2018/03/1521581382.jpg" class="entry-thumb" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521581382.jpg 942w, http://cronio.sv/wp-content/uploads/2018/03/1521581382-300x128.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/1521581382-768x328.jpg 768w" sizes="(max-width: 942px) 100vw, 942px" />						</a>
					</div>
					<div class="sa-meta-info-container">
						<div class="sa-meta-align">
							<div class="sa-big-grid-meta">
								<div class="svc_port_cat"><a>Internacionales</a></div>								<h3 class="entry-title sa-module-title"><a href="http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/">Mujer se opera los glúteos y ahora no puede sentarse</a></h3>
							</div>
						</div>
					</div>
				</div>
					
						<div class="sa-big-grid-post-1 sa-big-grid-post sa-small-thumb">
						<div class="svc_share">                            
		<i class="fa fa-share-alt"></i>
		<div class="svc_share-box full-color">
		  <ul class="s8-social">
			<li class="facebook">
				<a href="https://www.facebook.com/sharer/sharer.php?u=http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/" target="_blank" title="">
					<i class="fa fa-facebook"></i>
				</a>
			</li>
			<li class="google">
				<a href="https://plusone.google.com/share?url=http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/" target="_blank" title="">
					<i class="fa fa-google-plus"></i>
				</a>
			</li>
			<li class="twitter">
				<a href="https://twitter.com/intent/tweet?text=&amp;url=http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/" target="_blank" title="">
					<i class="fa fa-twitter"></i>
				</a>
			</li>
		  </ul>
		</div>
	</div>
						<div class="sa-module-thumb">
						<a href="http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/" target="_self">
							<img width="627" height="360" src="http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua.jpg" class="entry-thumb" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua.jpg 627w, http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua-300x172.jpg 300w" sizes="(max-width: 627px) 100vw, 627px" />						</a>
					</div>
					<div class="sa-meta-info-container">
						<div class="sa-meta-align">
							<div class="sa-big-grid-meta">
								<div class="svc_port_cat"><a>Judicial</a></div>								<h3 class="entry-title sa-module-title"><a href="http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/">Cámara ordena que se repita el juicio en el caso de la tregua entre pandillas</a></h3>
							</div>
						</div>
					</div>
				</div>
					
						<div class="sa-big-grid-post-1 sa-big-grid-post sa-small-thumb">
						<div class="svc_share">                            
		<i class="fa fa-share-alt"></i>
		<div class="svc_share-box full-color">
		  <ul class="s8-social">
			<li class="facebook">
				<a href="https://www.facebook.com/sharer/sharer.php?u=http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/" target="_blank" title="">
					<i class="fa fa-facebook"></i>
				</a>
			</li>
			<li class="google">
				<a href="https://plusone.google.com/share?url=http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/" target="_blank" title="">
					<i class="fa fa-google-plus"></i>
				</a>
			</li>
			<li class="twitter">
				<a href="https://twitter.com/intent/tweet?text=&amp;url=http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/" target="_blank" title="">
					<i class="fa fa-twitter"></i>
				</a>
			</li>
		  </ul>
		</div>
	</div>
						<div class="sa-module-thumb">
						<a href="http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/" target="_self">
							<img width="640" height="438" src="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438.jpg" class="entry-thumb" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438.jpg 640w, http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-300x205.jpg 300w" sizes="(max-width: 640px) 100vw, 640px" />						</a>
					</div>
					<div class="sa-meta-info-container">
						<div class="sa-meta-align">
							<div class="sa-big-grid-meta">
								<div class="svc_port_cat"><a>Internacionales</a></div>								<h3 class="entry-title sa-module-title"><a href="http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/">Empleado de zoológico muere tras ser atacado por un león</a></h3>
							</div>
						</div>
					</div>
				</div>
		</div>
				
				
				
				
				
				<div class="clearfix"></div>
		</div>
	</div>
	</div>
	<script>
	jQuery(document).ready(function(){		
		jQuery('#svc_post_grid_740').imagesLoaded( function() {
			jQuery('#svc_post_grid_list_container_740').show();
			jQuery('#svc_mask_740').hide();
			
		});
	});
</script>
		<div class="mvp-main-box">
		<section id="mvp-feat1-wrap" class="left relative">
			<div class="mvp-feat1-right-out left relative">
				<div class="mvp-feat1-right-in">
					<div class="mvp-feat1-main left relative">
						<div class="mvp-feat1-left-wrap relative">
															<a href="http://cronio.sv/nacionales/pnc-captura-14-pandilleros-ahuachapan/" rel="bookmark">
								<div class="mvp-feat1-feat-wrap left relative">
									<div class="mvp-feat1-feat-img left relative">
																					<img width="560" height="211" src="http://cronio.sv/wp-content/uploads/2018/03/DYw8zE_WAAAzl2R-560x211.jpg" class="attachment-mvp-port-thumb size-mvp-port-thumb wp-post-image" alt="" />																													</div><!--mvp-feat1-feat-img-->
									<div class="mvp-feat1-feat-text left relative">
										<div class="mvp-cat-date-wrap left relative">
											<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 7 horas</span>
										</div><!--mvp-cat-date-wrap-->
																					<h2 class="mvp-stand-title">PNC captura a 14 pandilleros en Ahuachapán </h2>
																				<p>Esta tarde de martes, autoridades de la Policía Nacional Civil (PNC) informaron sobre la captura de 10 criminales, la privación...</p>
									</div><!--mvp-feat1-feat-text-->
								</div><!--mvp-feat1-feat-wrap-->
								</a>
														<div class="mvp-feat1-sub-wrap left relative">
																	<a href="http://cronio.sv/nacionales/pnc-captura-medico-quien-acusado-abusar-una-joven-usulutan/" rel="bookmark">
									<div class="mvp-feat1-sub-cont left relative">
										<div class="mvp-feat1-sub-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/1521575580-590x354.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521575580-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/1521575580-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521575580-400x240.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521575580-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521575580-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-feat1-sub-img-->
										<div class="mvp-feat1-sub-text">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 9 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>PNC captura a Medico quien es acusado de abusar de una joven en Usulután</h2>
										</div><!--mvp-feat1-sub-text-->
									</div><!--mvp-feat1-sub-cont-->
									</a>
																	<a href="http://cronio.sv/nacionales/sucesos/hombre-cae-del-cuarto-piso-del-hospital-zacamil-del-isss/" rel="bookmark">
									<div class="mvp-feat1-sub-cont left relative">
										<div class="mvp-feat1-sub-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-590x354.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-400x240.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/2018032012183479734-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-feat1-sub-img-->
										<div class="mvp-feat1-sub-text">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Sucesos</span><span class="mvp-cd-date left relative">Hace 12 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Hombre cae del cuarto piso del hospital Zacamil del ISSS</h2>
										</div><!--mvp-feat1-sub-text-->
									</div><!--mvp-feat1-sub-cont-->
									</a>
															</div><!--mvp-feat1-sub-wrap-->
						</div><!--mvp-feat1-left-wrap-->
						<div class="mvp-feat1-mid-wrap left relative">
							<h3 class="mvp-feat1-pop-head"><span class="mvp-feat1-pop-head">Lo Más Leído</span></h3>
							<div class="mvp-feat1-pop-wrap left relative">
																	<a href="http://cronio.sv/nacionales/probidad-encuentra-indicios-enriquecimiento-ilicito-nayib-bukele-luis-mario-rodriguez-corte-plena-definir-juicios-este-martes/" rel="bookmark">
									<div class="mvp-feat1-pop-cont left relative">
																					<div class="mvp-feat1-pop-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/foto-ok-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/foto-ok-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/foto-ok-300x180.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/foto-ok-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/foto-ok.jpg 722w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/foto-ok-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/foto-ok-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/foto-ok-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																							</div><!--mvp-feat1-pop-img-->
																				<div class="mvp-feat1-pop-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Judicial</span><span class="mvp-cd-date left relative">Hace 2 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Probidad encuentra indicios de enriquecimiento ilícito contra Nayib Bukele y Luis Mario Rodríguez, Corte Plena por definir juicios este martes</h2>
										</div><!--mvp-feat1-pop-text-->
									</div><!--mvp-feat1-pop-cont-->
									</a>
																	<a href="http://cronio.sv/nacionales/matan-dueno-taller-automotriz-mejicanos/" rel="bookmark">
									<div class="mvp-feat1-pop-cont left relative">
																					<div class="mvp-feat1-pop-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/mejicanos-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/mejicanos-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/mejicanos-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/mejicanos-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/mejicanos-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/mejicanos-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																							</div><!--mvp-feat1-pop-img-->
																				<div class="mvp-feat1-pop-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 3 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Matan a dueño de taller automotriz en Mejicanos</h2>
										</div><!--mvp-feat1-pop-text-->
									</div><!--mvp-feat1-pop-cont-->
									</a>
																	<a href="http://cronio.sv/nacionales/ejecutan-dos-hombres-sonsonate/" rel="bookmark">
									<div class="mvp-feat1-pop-cont left relative">
																					<div class="mvp-feat1-pop-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/muertos-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/muertos-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/muertos-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/muertos-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/muertos-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/muertos-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																							</div><!--mvp-feat1-pop-img-->
																				<div class="mvp-feat1-pop-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 3 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Ejecutan a dos hombres en Sonsonate</h2>
										</div><!--mvp-feat1-pop-text-->
									</div><!--mvp-feat1-pop-cont-->
									</a>
																	<a href="http://cronio.sv/tendencias/jetset/ezequiel-garay-tamara-gorro-posan-desnudos-instagram/" rel="bookmark">
									<div class="mvp-feat1-pop-cont left relative">
																					<div class="mvp-feat1-pop-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																							</div><!--mvp-feat1-pop-img-->
																				<div class="mvp-feat1-pop-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 2 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Ezequiel Garay y Tamara Gorro posan desnudos para Instagram</h2>
										</div><!--mvp-feat1-pop-text-->
									</div><!--mvp-feat1-pop-cont-->
									</a>
																	<a href="http://cronio.sv/tendencias/jetset/revelan-foto-inedita-selena-quintanilla-luis-miguel/" rel="bookmark">
									<div class="mvp-feat1-pop-cont left relative">
																					<div class="mvp-feat1-pop-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																							</div><!--mvp-feat1-pop-img-->
																				<div class="mvp-feat1-pop-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 17 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Revelan foto inédita de Selena Quintanilla con Luis Miguel</h2>
										</div><!--mvp-feat1-pop-text-->
									</div><!--mvp-feat1-pop-cont-->
									</a>
															</div><!--mvp-feat1-pop-wrap-->
						</div><!--mvp-feat1-mid-wrap-->
					</div><!--mvp-feat1-main-->
				</div><!--mvp-feat1-right-in-->
				<div class="mvp-feat1-right-wrap left relative">

						<section id="mvp_flex_widget-3" class="mvp-side-widget mvp_flex_widget"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">CronioTV</span></h4></div>
		<div class="mvp-widget-flex-wrap left relative">
									<div class="mvp-flex-story-wrap left relative">
																																		<a href="http://cronio.sv/croniotv/alejandro-gutman-presidente-la-fundacion-forever-compartiendo-tema-la-cultura-la-integracion/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-col mvp-flex-col-noad">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/DYqUpCIVMAAv4JZ-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																													<div class="mvp-vid-box-wrap mvp-vid-marg">
																<i class="fa fa-2 fa-play" aria-hidden="true"></i>
															</div><!--mvp-vid-box-wrap-->
																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 2 días</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Alejandro Gutman, Presidente de la Fundación Forever, compartiendo el tema de la Cultura de la Integración</h2>
															<p>#ENVIVO EL SALVADOR TODAY con Alejandro Gutman, Presidente de la Fundación Forever, compartiendo el tema de la Cultura de la Integración....</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/croniotv/rodolfo-semsch-analista-experto-desarrollo-humano/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-col mvp-flex-col-noad">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/64c96a84-6227-4cc9-a7d7-97dd1a9dc68a-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																													<div class="mvp-vid-box-wrap mvp-vid-marg">
																<i class="fa fa-2 fa-play" aria-hidden="true"></i>
															</div><!--mvp-vid-box-wrap-->
																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 5 días</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Rodolfo Semsch, analista y experto en desarrollo humano</h2>
															<p>#ENVIVO EL SALVADOR TODAY con RODOLFO SEMSCH, ANALISTA Y EXPERTO EN DESARROLLO HUMANO. Envíe sus preguntas y comentarios a @croniosv o...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/croniotv/youtuberdad-diana-granadino-gerente-comercial-global-alimentos/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-col mvp-flex-col-noad">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/DYWH76iV4AA8S_y-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																													<div class="mvp-vid-box-wrap mvp-vid-marg">
																<i class="fa fa-2 fa-play" aria-hidden="true"></i>
															</div><!--mvp-vid-box-wrap-->
																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 6 días</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">YOUTUBERDAD con Diana Granadino, Gerente Relaciones Corporativas de Global Alimentos</h2>
															<p>#ENVIVO YOUTUBERDAD con Diana Granadino, Gerente comercial de Global Alimentos. Escríbanos a @croniosv o llámenos al Cronio WhatsApp 7017-4887. DANOS LIKE,...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																														</div><!--mvp-flex-story-wrap-->
					</div><!--mvp-widget-flex-wrap-->

		</section>
											<div class="mvp-feat1-list-ad left relative">
							<span class="mvp-ad-label">Advertisements</span>
							<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 300x250 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:300px;height:250px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="4286918273"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>						</div><!--mvp-feat1-list-ad-->
					

					

						

				</div><!--mvp-feat1-right-wrap-->
			</div><!--mvp-feat1-right-out-->
		</section><!--mvp-feat1-wrap-->
	</div><!--mvp-main-box-->
	<div id="mvp-home-widget-wrap" class="left relative">
					<section id="mvp_home_feat2_widget-2" class="mvp-widget-home left relative mvp_home_feat2_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Nacionales</span></h4></div>
			<div class="mvp-widget-feat2-wrap left relative">
				<div class="mvp-widget-feat2-out left relative">
					<div class="mvp-widget-feat2-in">
						<div class="mvp-widget-feat2-main left relative">
															<div class="mvp-widget-feat2-left left relative mvp-widget-feat2-left-alt">
																																													<a href="http://cronio.sv/nacionales/judicial/investigadores-la-pnc-capturados-matar-agente-alterar-la-escena-del-crimen/" rel="bookmark">
											<div class="mvp-widget-feat2-left-cont left relative">
												<div class="mvp-feat1-feat-img left relative">
																											<img width="560" height="541" src="http://cronio.sv/wp-content/uploads/2018/03/esposados-560x541.jpg" class="attachment-mvp-port-thumb size-mvp-port-thumb wp-post-image" alt="" />																																						</div><!--mvp-feat1-feat-img-->
												<div class="mvp-feat1-feat-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">Judicial</span><span class="mvp-cd-date left relative">Hace 7 horas</span>
													</div><!--mvp-cat-date-wrap-->
																											<h2 class="mvp-stand-title">Investigadores de la PNC son capturados por matar a otro agente y alterar la escena del crimen</h2>
																										<p>Dos elementos de la Unidad de Investigaciones de la Policía Nacional Civil (PNC), identificados como José Durán y David Barahona...</p>
												</div><!--mvp-feat1-feat-text-->
											</div><!--mvp-widget-feat2-left-cont-->
											</a>
																																		</div><!--mvp-widget-feat2-left-->
							<div class="mvp-widget-feat2-right left relative">
																											<a href="http://cronio.sv/nacionales/judicial/juez-ordena-jorge-hernandez-conciliara-periodistas-quienes-habria-retenido-cuotas-seguro-social-afp/" rel="bookmark">
										<div class="mvp-widget-feat2-right-cont left relative">
											<div class="mvp-widget-feat2-right-img left relative">
																									<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />													<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/Jorge-hernández-7-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																			</div><!--mvp-widget-feat2-right-img-->
											<div class="mvp-widget-feat2-right-text left relative">
												<div class="mvp-cat-date-wrap left relative">
													<span class="mvp-cd-cat left relative">Judicial</span><span class="mvp-cd-date left relative">Hace 8 horas</span>
												</div><!--mvp-cat-date-wrap-->
												<h2>Juez ordena que Jorge Hernández, conciliara con algunos periodistas a quienes habría retenido cuotas de Seguro Social y AFP</h2>
											</div><!--mvp-widget-feat2-right-text-->
										</div><!--mvp-widget-feat2-right-cont-->
										</a>
																			<a href="http://cronio.sv/nacionales/bulevar-venezuela-cerrado-accidente-transito/" rel="bookmark">
										<div class="mvp-widget-feat2-right-cont left relative">
											<div class="mvp-widget-feat2-right-img left relative">
																									<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521586878-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521586878-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521586878-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />													<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/1521586878-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521586878-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/1521586878-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																			</div><!--mvp-widget-feat2-right-img-->
											<div class="mvp-widget-feat2-right-text left relative">
												<div class="mvp-cat-date-wrap left relative">
													<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 8 horas</span>
												</div><!--mvp-cat-date-wrap-->
												<h2>Bulevar Venezuela cerrado por accidente de tránsito</h2>
											</div><!--mvp-widget-feat2-right-text-->
										</div><!--mvp-widget-feat2-right-cont-->
										</a>
																								</div><!--mvp-widget-feat2-right-->
						</div><!--mvp-widget-feat2-main-->
					</div><!--mvp-widget-feat2-in-->
					<div class="mvp-widget-feat2-side left relative">
													<div class="mvp-widget-feat2-side-ad left relative">
								<span class="mvp-ad-label">Advertisement</span>
								<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 300x250 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:300px;height:250px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="4286918273"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>							</div><!--mvp-widget-feat2-side-ad-->
												<div class="mvp-widget-feat2-side-list left relative">
							<div class="mvp-feat1-list left relative">
																											<a href="http://cronio.sv/nacionales/judicial/camara-ordena-se-repita-juicio-caso-la-tregua-pandillas/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua-80x80.jpg" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/Audiencia-caso-tregua-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Judicial</span><span class="mvp-cd-date left relative">Hace 10 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Cámara ordena que se repita el juicio en el caso de la tregua entre pandillas</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																			<a href="http://cronio.sv/nacionales/sujetos-capturados-compartir-material-intimo-redes-sociales/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/capturados-80x80.jpg" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/capturados-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/capturados-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 11 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Sujetos son capturados por compartir material intimo en redes sociales</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																			<a href="http://cronio.sv/nacionales/menor-edad-herido-bala-disputa-comerciantes-agentes-del-cam-santa-tecla/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/IMG-20180320-WA0015-300x169-1-80x80.jpg" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/IMG-20180320-WA0015-300x169-1-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/IMG-20180320-WA0015-300x169-1-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Nacionales</span><span class="mvp-cd-date left relative">Hace 12 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Menor de edad es herido de bala en disputa entre comerciantes y agentes del CAM en Santa Tecla</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																								</div><!--mvp-feat1-list-->
															<a href="http://cronio.sv/category/nacionales/">
								<div class="mvp-widget-feat2-side-more-but left relative">
									<span class="mvp-widget-feat2-side-more">More Nacionales</span><i class="fa fa-long-arrow-right" aria-hidden="true"></i>
								</div><!--mvp-widget-feat2-side-more-but-->
								</a>
													</div><!--mvp-widget-feat2-side-list-->
					</div><!--mvp-widget-feat2-side-->
				</div><!--mvp-widget-feat2-out-->
			</div><!--mvp-widget-feat2-wrap-->

		</div></section><section id="mvp_ad_widget-8" class="mvp-widget-home left relative mvp_ad_widget"><div class="mvp-main-box">			<div class="mvp-widget-ad left relative">
				<span class="mvp-ad-label">Advertisement</span>
				<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 728*90 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:728px;height:90px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="6030835660"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>			</div><!--mvp-widget-ad-->
		</div></section>
	<section class="mvp-widget-home left relative">
		<div class="mvp-widget-dark-wrap left relative">
			<div class="mvp-main-box">
				<div class="mvp-widget-home-head">
					<h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">CronioTV</span></h4>
				</div><!--mvp-widget-home-head-->
				<div class="mvp-widget-dark-main left relative">
					<div class="mvp-widget-dark-left left relative">
																														<a href="http://cronio.sv/croniotv/christian-aparicio-docente-universitario-habla-del-marketing-politico-pais/" rel="bookmark">
									<div class="mvp-widget-dark-feat left relative">
										<div class="mvp-widget-dark-feat-img left relative">
																							<img width="739" height="327" src="http://cronio.sv/wp-content/uploads/2018/03/e74e20c2-8651-4e96-9561-c94bd26851de.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/e74e20c2-8651-4e96-9561-c94bd26851de.jpg 739w, http://cronio.sv/wp-content/uploads/2018/03/e74e20c2-8651-4e96-9561-c94bd26851de-300x133.jpg 300w" sizes="(max-width: 739px) 100vw, 739px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/e74e20c2-8651-4e96-9561-c94bd26851de-400x240.jpg" class="mvp-mob-img lazy wp-post-image" alt="" />																																		<div class="mvp-vid-box-wrap mvp-vid-marg">
													<i class="fa fa-2 fa-play" aria-hidden="true"></i>
												</div><!--mvp-vid-box-wrap-->
																					</div><!--mvp-widget-dark-feat-img-->
										<div class="mvp-widget-dark-feat-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 7 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Christian Aparicio, docente universitario habla del marketing político en el país</h2>
										</div><!--mvp-widget-dark-feat-text-->
									</div><!--mvp-widget-dark-feat-->
									</a>
																										</div><!--mvp-widget-dark-left-->
					<div class="mvp-widget-dark-right left relative">
																					<a href="http://cronio.sv/croniotv/envivo-nuevo-episodio-cronio-al-extremo-josue-herrera/" rel="bookmark">
								<div class="mvp-widget-dark-sub left relative">
																			<div class="mvp-widget-dark-sub-out right relative">
											<div class="mvp-widget-dark-sub-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-150x150.jpg 150w, http://cronio.sv/wp-content/uploads/2018/03/29101444_1476336562494407_2574071061242970112_n-560x556.jpg 560w" sizes="(max-width: 80px) 100vw, 80px" />																									<div class="mvp-vid-box-wrap mvp-vid-box-small mvp-vid-marg-small">
														<i class="fa fa-2 fa-play" aria-hidden="true"></i>
													</div><!--mvp-vid-box-wrap-->
																							</div><!--mvp-widget-dark-sub-img-->
											<div class="mvp-widget-dark-sub-in">
												<div class="mvp-widget-dark-sub-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 1 semana</span>
													</div><!--mvp-cat-date-wrap-->
													<h2>#ENVIVO Un nuevo episodio de Cronio al Extremo, con Josué Herrera</h2>
												</div><!--mvp-widget-dark-sub-text-->
											</div><!--mvp-widget-dark-sub-in-->
										</div><!--mvp-widget-dark-sub-out-->
																	</div><!--mvp-widget-dark-sub-->
								</a>
															<a href="http://cronio.sv/croniotv/felix-ulloa-exmagistrado-analista-politico-habla-del-acontecer-politico-tras-las-elecciones-2018/" rel="bookmark">
								<div class="mvp-widget-dark-sub left relative">
																			<div class="mvp-widget-dark-sub-out right relative">
											<div class="mvp-widget-dark-sub-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/2b943b3f-8ab0-425f-b911-743d1de4a25f-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																									<div class="mvp-vid-box-wrap mvp-vid-box-small mvp-vid-marg-small">
														<i class="fa fa-2 fa-play" aria-hidden="true"></i>
													</div><!--mvp-vid-box-wrap-->
																							</div><!--mvp-widget-dark-sub-img-->
											<div class="mvp-widget-dark-sub-in">
												<div class="mvp-widget-dark-sub-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 1 semana</span>
													</div><!--mvp-cat-date-wrap-->
													<h2>Félix Ulloa, exmagistrado y analista político habla del acontecer político tras las elecciones 2018</h2>
												</div><!--mvp-widget-dark-sub-text-->
											</div><!--mvp-widget-dark-sub-in-->
										</div><!--mvp-widget-dark-sub-out-->
																	</div><!--mvp-widget-dark-sub-->
								</a>
															<a href="http://cronio.sv/uncategorized/eduardo-escobar-isd-analizando-los-datos-preliminares-la-eleccion-legislativa-municipal/" rel="bookmark">
								<div class="mvp-widget-dark-sub left relative">
																			<div class="mvp-widget-dark-sub-out right relative">
											<div class="mvp-widget-dark-sub-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Captura-6-400x240.png" class="mvp-reg-img lazy wp-post-image" alt="" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Captura-6-80x80.png" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Captura-6-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/Captura-6-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />																									<div class="mvp-vid-box-wrap mvp-vid-box-small mvp-vid-marg-small">
														<i class="fa fa-2 fa-play" aria-hidden="true"></i>
													</div><!--mvp-vid-box-wrap-->
																							</div><!--mvp-widget-dark-sub-img-->
											<div class="mvp-widget-dark-sub-in">
												<div class="mvp-widget-dark-sub-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">CronioTV</span><span class="mvp-cd-date left relative">Hace 2 semanas</span>
													</div><!--mvp-cat-date-wrap-->
													<h2>Eduardo Escobar, de Acción Ciudadana, analizando los datos preliminares de la Elección Legislativa y Municipal</h2>
												</div><!--mvp-widget-dark-sub-text-->
											</div><!--mvp-widget-dark-sub-in-->
										</div><!--mvp-widget-dark-sub-out-->
																	</div><!--mvp-widget-dark-sub-->
								</a>
															<a href="http://cronio.sv/uncategorized/elecciones-legislativas-municipales-salvador-2/" rel="bookmark">
								<div class="mvp-widget-dark-sub left relative">
																			<div class="mvp-widget-dark-sub-out right relative">
											<div class="mvp-widget-dark-sub-img left relative">
												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/programa-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/programa-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/programa-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/programa-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																									<div class="mvp-vid-box-wrap mvp-vid-box-small mvp-vid-marg-small">
														<i class="fa fa-2 fa-play" aria-hidden="true"></i>
													</div><!--mvp-vid-box-wrap-->
																							</div><!--mvp-widget-dark-sub-img-->
											<div class="mvp-widget-dark-sub-in">
												<div class="mvp-widget-dark-sub-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">Uncategorized</span><span class="mvp-cd-date left relative">Hace 2 semanas</span>
													</div><!--mvp-cat-date-wrap-->
													<h2>ELECCIONES LEGISLATIVAS Y MUNICIPALES DE EL SALVADOR</h2>
												</div><!--mvp-widget-dark-sub-text-->
											</div><!--mvp-widget-dark-sub-in-->
										</div><!--mvp-widget-dark-sub-out-->
																	</div><!--mvp-widget-dark-sub-->
								</a>
																		</div><!--mvp-widget-dark-right-->
				</div><!--mvp-widget-dark-main-->
			</div><!--mvp-main-box-->
		</div><!--mvp-widget-dark-wrap-->
	</section><!--mvp-widget-home-->

		<section id="mvp_ad_widget-5" class="mvp-widget-home left relative mvp_ad_widget"><div class="mvp-main-box">			<div class="mvp-widget-ad left relative">
				<span class="mvp-ad-label">Advertisement</span>
				<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 728*90 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:728px;height:90px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="6030835660"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>			</div><!--mvp-widget-ad-->
		</div></section><section id="mvp_home_feat1_widget-2" class="mvp-widget-home left relative mvp_home_feat1_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Política</span></h4></div>
			<div class="mvp-widget-feat1-wrap left relative">
									<div class="mvp-widget-feat1-cont left relative">
																														<a href="http://cronio.sv/politica/carlos-caceres-anuncia-sera-nuevo-embajador-mexico/" rel="bookmark">
									<div class="mvp-widget-feat1-top-story left relative">
										<div class="mvp-widget-feat1-top-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-590x354.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-400x240.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/Ministro_Hacienda-Carlos_Cáceres-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-widget-feat1-top-img-->
										<div class="mvp-widget-feat1-top-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 7 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Carlos Cáceres, anuncia que sera el nuevo Embajador en México</h2>
										</div><!--mvp-widget-feat1-top-text-->
									</div><!--mvp-widget-feat1-top-story-->
									</a>
																	<a href="http://cronio.sv/politica/lopez-davidson-cambios-gobierno-fue-reciclaje-decorativo-los-mismos-funcionarios/" rel="bookmark">
									<div class="mvp-widget-feat1-top-story left relative">
										<div class="mvp-widget-feat1-top-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/tavo-590x354.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tavo-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/tavo-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tavo-400x240.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tavo-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/tavo-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-widget-feat1-top-img-->
										<div class="mvp-widget-feat1-top-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 10 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>López Davidson: &#8220;Cambios en el Gobierno fue un reciclaje decorativo de los mismos funcionarios&#8221;</h2>
										</div><!--mvp-widget-feat1-top-text-->
									</div><!--mvp-widget-feat1-top-story-->
									</a>
																										</div><!--mvp-widget-feat1-cont-->
													<div class="mvp-widget-feat1-cont left relative">
																														<a href="http://cronio.sv/politica/smartmatic-sera-demanda-tse-confirma-julio-olivo/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/tseconferencia-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 15 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Smartmatic será demanda por el TSE confirma Julio Olivo</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/politica/ya-no-habran-mas-cambios-gabinete-gobierno-dice-roberto-lorenzana/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/LORENZANA-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 16 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Ya no habrán más cambios en el gabinete de gobierno dice Roberto Lorenzana</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/politica/norman-quijano-aspira-la-presidencia-la-asamblea-legislativa-gracias-al-voto-popular/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/Norman-Quijano-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 1 día</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Norman Quijano aspira a la presidencia de la Asamblea Legislativa gracias al voto popular</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/politica/eugenio-chicas-tras-destituido-cargo-no-pudimos-bien-trabajo-comunicar-las-acciones-del-gobierno/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-400x240.png" class="mvp-reg-img lazy wp-post-image" alt="Eugenio Chicas tras ser destituido de su cargo: No pudimos hacer bien nuestro trabajo de comunicar las acciones del Gobierno" srcset="http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-400x240.png 400w, http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-1000x600.png 1000w, http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-590x354.png 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-80x80.png" class="mvp-mob-img lazy wp-post-image" alt="Eugenio Chicas tras ser destituido de su cargo: No pudimos hacer bien nuestro trabajo de comunicar las acciones del Gobierno" srcset="http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/Eugenio-Chicas-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Política</span><span class="mvp-cd-date left relative">Hace 1 día</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Eugenio Chicas tras ser destituido de su cargo: No pudimos hacer bien nuestro trabajo de comunicar las acciones del Gobierno</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																										</div><!--mvp-widget-feat1-cont-->
							</div><!--mvp-widget-feat1-wrap-->

		</div></section><section id="mvp_ad_widget-6" class="mvp-widget-home left relative mvp_ad_widget"><div class="mvp-main-box">			<div class="mvp-widget-ad left relative">
				<span class="mvp-ad-label">Advertisement</span>
				<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 728*90 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:728px;height:90px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="6030835660"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>			</div><!--mvp-widget-ad-->
		</div></section><section id="mvp_home_feat2_widget-3" class="mvp-widget-home left relative mvp_home_feat2_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Internacionales</span></h4></div>
			<div class="mvp-widget-feat2-wrap left relative">
				<div class="mvp-widget-feat2-out left relative">
					<div class="mvp-widget-feat2-in">
						<div class="mvp-widget-feat2-main left relative">
															<div class="mvp-widget-feat2-left left relative">
																																													<a href="http://cronio.sv/internacionales/pareja-sorprendida-azafata-tenian-intimidad-avion/" rel="bookmark">
											<div class="mvp-widget-feat2-left-cont left relative">
												<div class="mvp-feat1-feat-img left relative">
																											<img width="560" height="375" src="http://cronio.sv/wp-content/uploads/2018/03/1521572499-560x375.jpg" class="attachment-mvp-port-thumb size-mvp-port-thumb wp-post-image" alt="" />																																						</div><!--mvp-feat1-feat-img-->
												<div class="mvp-feat1-feat-text left relative">
													<div class="mvp-cat-date-wrap left relative">
														<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 7 horas</span>
													</div><!--mvp-cat-date-wrap-->
																											<h2 class="mvp-stand-title">Pareja es sorprendida por azafata mientras tenían intimidad en un avión</h2>
																										<p>Durante un viaje aéreo hacia México la empleada de una aerolínea Entró al baño y encontró a un hombre y...</p>
												</div><!--mvp-feat1-feat-text-->
											</div><!--mvp-widget-feat2-left-cont-->
											</a>
																																		</div><!--mvp-widget-feat2-left-->
							<div class="mvp-widget-feat2-right left relative">
																											<a href="http://cronio.sv/internacionales/mujer-se-opera-los-gluteos-ahora-no-puede-sentarse/" rel="bookmark">
										<div class="mvp-widget-feat2-right-cont left relative">
											<div class="mvp-widget-feat2-right-img left relative">
																									<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521581382-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521581382-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521581382-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />													<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/1521581382-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521581382-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/1521581382-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																			</div><!--mvp-widget-feat2-right-img-->
											<div class="mvp-widget-feat2-right-text left relative">
												<div class="mvp-cat-date-wrap left relative">
													<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 9 horas</span>
												</div><!--mvp-cat-date-wrap-->
												<h2>Mujer se opera los glúteos y ahora no puede sentarse</h2>
											</div><!--mvp-widget-feat2-right-text-->
										</div><!--mvp-widget-feat2-right-cont-->
										</a>
																			<a href="http://cronio.sv/internacionales/empleado-zoologico-muere-tras-atacado-leon/" rel="bookmark">
										<div class="mvp-widget-feat2-right-cont left relative">
											<div class="mvp-widget-feat2-right-img left relative">
																									<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />													<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/lo-640x438-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																			</div><!--mvp-widget-feat2-right-img-->
											<div class="mvp-widget-feat2-right-text left relative">
												<div class="mvp-cat-date-wrap left relative">
													<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 11 horas</span>
												</div><!--mvp-cat-date-wrap-->
												<h2>Empleado de zoológico muere tras ser atacado por un león</h2>
											</div><!--mvp-widget-feat2-right-text-->
										</div><!--mvp-widget-feat2-right-cont-->
										</a>
																								</div><!--mvp-widget-feat2-right-->
						</div><!--mvp-widget-feat2-main-->
					</div><!--mvp-widget-feat2-in-->
					<div class="mvp-widget-feat2-side left relative">
													<div class="mvp-widget-feat2-side-ad left relative">
								<span class="mvp-ad-label">Advertisement</span>
								<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 300x250 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:300px;height:250px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="4286918273"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>							</div><!--mvp-widget-feat2-side-ad-->
												<div class="mvp-widget-feat2-side-list left relative">
							<div class="mvp-feat1-list left relative">
																											<a href="http://cronio.sv/internacionales/hombre-paso-25-anos-corredor-la-muerte-tras-condenado-pruebas-falsas-abusar-asesinar-una-bebe/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/cdn1.uvnimg-80x80.png" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/cdn1.uvnimg-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/cdn1.uvnimg-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 12 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Hombre pasó 25 años en el corredor de la muerte tras ser condenado con pruebas falsas de abusar y asesinar a una bebé</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																			<a href="http://cronio.sv/internacionales/nicolas-sarkozy-detenido-la-presunta-financiacion-ilegal-campana-2007/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/imagen-sin-titulo-80x80.jpg" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/imagen-sin-titulo-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/imagen-sin-titulo-150x150.jpg 150w, http://cronio.sv/wp-content/uploads/2018/03/imagen-sin-titulo-560x560.jpg 560w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 19 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Nicolás Sarkozy, detenido por la presunta financiación ilegal de su campaña en 2007</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																			<a href="http://cronio.sv/internacionales/investigan-tiroteo-una-escuela-secundaria-maryland/" rel="bookmark">
										<div class="mvp-feat1-list-cont left relative">
																							<div class="mvp-feat1-list-out relative">
													<div class="mvp-feat1-list-img left relative">
														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/DYu-x_xW4AE8U25-80x80.jpg" class="attachment-mvp-small-thumb size-mvp-small-thumb wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/DYu-x_xW4AE8U25-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/DYu-x_xW4AE8U25-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />													</div><!--mvp-feat1-list-img-->
													<div class="mvp-feat1-list-in">
														<div class="mvp-feat1-list-text">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Internacionales</span><span class="mvp-cd-date left relative">Hace 19 horas</span>
															</div><!--mvp-cat-date-wrap-->
															<h2>Investigan un tiroteo en una escuela secundaria en Maryland</h2>
														</div><!--mvp-feat1-list-text-->
													</div><!--mvp-feat1-list-in-->
												</div><!--mvp-feat1-list-out-->
																					</div><!--mvp-feat1-list-cont-->
										</a>
																								</div><!--mvp-feat1-list-->
															<a href="http://cronio.sv/category/internacionales/">
								<div class="mvp-widget-feat2-side-more-but left relative">
									<span class="mvp-widget-feat2-side-more">More Internacionales</span><i class="fa fa-long-arrow-right" aria-hidden="true"></i>
								</div><!--mvp-widget-feat2-side-more-but-->
								</a>
													</div><!--mvp-widget-feat2-side-list-->
					</div><!--mvp-widget-feat2-side-->
				</div><!--mvp-widget-feat2-out-->
			</div><!--mvp-widget-feat2-wrap-->

		</div></section><section id="mvp_home_feat1_widget-3" class="mvp-widget-home left relative mvp_home_feat1_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Deportes</span></h4></div>
			<div class="mvp-widget-feat1-wrap left relative">
									<div class="mvp-widget-feat1-cont left relative">
																														<a href="http://cronio.sv/deportes/internacionales-deportes/messi-luce-la-nueva-indumentaria-alternativa-argentina-mundial-rusia-2018/" rel="bookmark">
									<div class="mvp-widget-feat1-top-story left relative">
										<div class="mvp-widget-feat1-top-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-590x354.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-400x240.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/ae3a7f2e-c7d9-4e7c-91f3-9368710f52a8_749_499-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-widget-feat1-top-img-->
										<div class="mvp-widget-feat1-top-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Internacionales -deportes</span><span class="mvp-cd-date left relative">Hace 13 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Messi luce la nueva indumentaria alternativa de Argentina para el Mundial Rusia 2018</h2>
										</div><!--mvp-widget-feat1-top-text-->
									</div><!--mvp-widget-feat1-top-story-->
									</a>
																	<a href="http://cronio.sv/deportes/internacionales-deportes/cristiano-ronaldo-no-nadie-mejor/" rel="bookmark">
									<div class="mvp-widget-feat1-top-story left relative">
										<div class="mvp-widget-feat1-top-img left relative">
																							<img width="590" height="354" src="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-590x354.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-400x240.jpg 400w" sizes="(max-width: 590px) 100vw, 590px" />												<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-400x240.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/hi-res-ff56c8d386e897e0bd3f71edf145900c_crop_north-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />																																</div><!--mvp-widget-feat1-top-img-->
										<div class="mvp-widget-feat1-top-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Internacionales -deportes</span><span class="mvp-cd-date left relative">Hace 18 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Cristiano Ronaldo: “No hay nadie mejor que yo”</h2>
										</div><!--mvp-widget-feat1-top-text-->
									</div><!--mvp-widget-feat1-top-story-->
									</a>
																										</div><!--mvp-widget-feat1-cont-->
													<div class="mvp-widget-feat1-cont left relative">
																														<a href="http://cronio.sv/deportes/real-madrid-arrolla-al-girona-6-3/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/madrid-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/madrid-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/madrid-300x180.jpg 300w, http://cronio.sv/wp-content/uploads/2018/03/madrid-590x354.jpg 590w, http://cronio.sv/wp-content/uploads/2018/03/madrid.jpg 700w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/madrid-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/madrid-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/madrid-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Deportes</span><span class="mvp-cd-date left relative">Hace 2 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>El Real Madrid arrolla al Girona 6-3</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/deportes/barca-se-impone-2-0-al-athletic-avanza-la-liga/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/barca-1-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/barca-1-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/barca-1-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/barca-1-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/barca-1-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/barca-1-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Deportes</span><span class="mvp-cd-date left relative">Hace 3 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>El Barca se impone 2-0 al Athletic y avanza en la Liga</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/deportes/messi-baila-celebrar-gol-frente-al-athletic/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/messi-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/messi-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/messi-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/messi-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/messi-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/messi-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/messi-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Deportes</span><span class="mvp-cd-date left relative">Hace 3 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>VIDEO Messi baila para celebrar su gol frente al Athletic</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/deportes/internacionales-deportes/neymar-jr-la-lesion-posible-boda-bruna-marquezine/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Neymar-400x240.png" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Neymar-400x240.png 400w, http://cronio.sv/wp-content/uploads/2018/03/Neymar-590x354.png 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Neymar-80x80.png" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Neymar-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/Neymar-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Internacionales -deportes</span><span class="mvp-cd-date left relative">Hace 5 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Neymar Jr. entre la lesión y su posible boda con Bruna Marquezine</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																										</div><!--mvp-widget-feat1-cont-->
							</div><!--mvp-widget-feat1-wrap-->

		</div></section><section id="mvp_ad_widget-7" class="mvp-widget-home left relative mvp_ad_widget"><div class="mvp-main-box">			<div class="mvp-widget-ad left relative">
				<span class="mvp-ad-label">Advertisement</span>
				<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 728*90 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:728px;height:90px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="6030835660"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>			</div><!--mvp-widget-ad-->
		</div></section><section id="mvp_home_feat1_widget-4" class="mvp-widget-home left relative mvp_home_feat1_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Tendencias</span></h4></div>
			<div class="mvp-widget-feat1-wrap left relative">
													<div class="mvp-widget-feat1-cont left relative">
																														<a href="http://cronio.sv/tendencias/jetset/will-smith-se-roba-show-al-ritmo-x-nick-jam-j-balvin/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Captura-20-400x240.png" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Captura-20-400x240.png 400w, http://cronio.sv/wp-content/uploads/2018/03/Captura-20-590x354.png 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Captura-20-80x80.png" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Captura-20-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/Captura-20-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 16 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>VIDEO: Will Smith se roba el show al ritmo de ´X´ de Nick Jam y J Balvin</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/tendencias/jetset/revelan-foto-inedita-selena-quintanilla-luis-miguel/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-1000x600.jpg 1000w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/5aaeb0d4efa06-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 17 horas</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Revelan foto inédita de Selena Quintanilla con Luis Miguel</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/tendencias/jetset/amaia-montero-exvocalista-la-oreja-van-gogh-luce-nuevo-rostro/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/amaia-montero-cambio-kDXF-U501316079844yLG-624x385@El-Comercio-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 1 día</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Amaia Montero, exvocalista de La Oreja de Van Gogh luce nuevo rostro</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																	<a href="http://cronio.sv/tendencias/jetset/ezequiel-garay-tamara-gorro-posan-desnudos-instagram/" rel="bookmark">
									<div class="mvp-widget-feat1-bot-story left relative">
										<div class="mvp-widget-feat1-bot-img left relative">
																							<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-400x240.jpg" class="mvp-reg-img lazy wp-post-image" alt="" />												<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-80x80.jpg" class="mvp-mob-img lazy wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/tamara-gorro-ezequiel-presenta-hijo-antonio-01_galeria_landscape-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																																</div><!--mvp-widget-feat1-bot-img-->
										<div class="mvp-widget-feat1-bot-text left relative">
											<div class="mvp-cat-date-wrap left relative">
												<span class="mvp-cd-cat left relative">Jetset</span><span class="mvp-cd-date left relative">Hace 2 días</span>
											</div><!--mvp-cat-date-wrap-->
											<h2>Ezequiel Garay y Tamara Gorro posan desnudos para Instagram</h2>
										</div><!--mvp-widget-feat1-bot-text-->
									</div><!--mvp-widget-feat1-bot-story-->
									</a>
																										</div><!--mvp-widget-feat1-cont-->
							</div><!--mvp-widget-feat1-wrap-->

		</div></section><section id="mvp_flex_widget-4" class="mvp-widget-home left relative mvp_flex_widget"><div class="mvp-main-box"><div class="mvp-widget-home-head"><h4 class="mvp-widget-home-title"><span class="mvp-widget-home-title">Redes</span></h4></div>
		<div class="mvp-widget-flex-wrap left relative">
							<div class="mvp-flex-side-out left relative">
					<div class="mvp-flex-side-in">
						<div class="mvp-flex-story-wrap left relative">
																																		<a href="http://cronio.sv/redes/viral-video-mono-desnuda-una-joven-turista/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1521478354-400x240.jpg" class="mvp-reg-img wp-post-image" alt="Mono desnuda a una joven turista" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521478354-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/1521478354-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/1521478354-80x80.jpg" class="mvp-mob-img wp-post-image" alt="Mono desnuda a una joven turista" srcset="http://cronio.sv/wp-content/uploads/2018/03/1521478354-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/1521478354-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Redes</span><span class="mvp-cd-date left relative">Hace 1 día</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">#VIRAL #VIDEO: Mono desnuda a una joven turista</h2>
															<p>Una incómoda situación, aunque ella se lo tomó con bastante humor, vivió una joven turista estadounidense mientras visitaba una localidad...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/redes/guatemala-captan-video-cuando-trabajador-bus-golpea-pasajera/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/Guatemala-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/Guatemala-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/Guatemala-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/Guatemala-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Redes</span><span class="mvp-cd-date left relative">Hace 3 días</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Guatemala: Captan en video cuando trabajador de bus que golpea a pasajera</h2>
															<p>Una mujer recibió un golpe de parte de un cobrador de bus porque se negó a pagar una parte del...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/redes/virales/mujer-da-luz-mar-rojo-impresionante-sucede/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/58-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/58-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/58-590x354.jpg 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/58-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/58-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/58-150x150.jpg 150w, http://cronio.sv/wp-content/uploads/2018/03/58-560x567.jpg 560w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Virales</span><span class="mvp-cd-date left relative">Hace 4 días</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Mujer da a luz en el mar rojo y esto impresionante sucede</h2>
															<p>Las imágenes de una turista rusa dando a luz en una playa de Dahab, en el mar Rojo (Egipto), se...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/redes/virales/sujeto-golpea-una-mujer-sin-conocerla-plena-via-publica/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/1520873216-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/1520873216-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/1520873216-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/1520873216-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Virales</span><span class="mvp-cd-date left relative">Hace 1 semana</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Sujeto golpea a una mujer sin conocerla en plena vía pública</h2>
															<p>En las últimas horas se ha vuelto viral un video que muestra el momento en que un hombre desconocido dio...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/redes/joven-ofrece-redes-sociales-relaciones-se-llevo-la-sorpresa-vida/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/65401-400x240.png" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/65401-400x240.png 400w, http://cronio.sv/wp-content/uploads/2018/03/65401-590x354.png 590w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/65401-80x80.png" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/65401-80x80.png 80w, http://cronio.sv/wp-content/uploads/2018/03/65401-150x150.png 150w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Redes</span><span class="mvp-cd-date left relative">Hace 1 semana</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Joven ofrece en redes sociales tener &#8220;relaciones&#8221; y se llevo la sorpresa de su vida</h2>
															<p>Qianjin Yeye, una joven china de 19 años de edad, se convirtió en estrella de internet por un día después...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																			<a href="http://cronio.sv/redes/virales/cientificos-captan-extrano-familiar-sonido-las-entranas-glaciar-antartico/" rel="bookmark">
																					<div class="mvp-flex-story left relative mvp-flex-row">
																																	<div class="mvp-flex-story-out right relative">
													<div class="mvp-flex-story-img left relative">
														<img width="400" height="240" src="http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-400x240.jpg" class="mvp-reg-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-400x240.jpg 400w, http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-560x338.jpg 560w" sizes="(max-width: 400px) 100vw, 400px" />														<img width="80" height="80" src="http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-80x80.jpg" class="mvp-mob-img wp-post-image" alt="" srcset="http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-80x80.jpg 80w, http://cronio.sv/wp-content/uploads/2018/03/650354-600-338-150x150.jpg 150w" sizes="(max-width: 80px) 100vw, 80px" />																											</div><!--mvp-flex-story-img--->
													<div class="mvp-flex-story-in">
														<div class="mvp-flex-story-text left relative">
															<div class="mvp-cat-date-wrap left relative">
																<span class="mvp-cd-cat left relative">Virales</span><span class="mvp-cd-date left relative">Hace 1 semana</span>
															</div><!--mvp-cat-date-wrap-->
															<h2 class="mvp-stand-title">Científicos captan un extraño (y familiar) sonido en las entrañas de un glaciar antártico</h2>
															<p>Un glaciólogo de un laboratorio de la Universidad de Rochester, Peter Neff ha publicado en su cuenta Twitter un video...</p>
														</div><!--mvp-flex-story-text--->
													</div><!--mvp-flex-story-in-->
												</div><!--mvp-flex-story-out-->
																					</div><!--mvp-flex-story-->
										</a>
																														</div><!--mvp-flex-story-wrap-->
					</div><!--mvp-flex-side-in-->
					<div class="mvp-flex-side-wrap left relative">
						<div class="mvp-flex-ad left relative">
							<span class="mvp-ad-label">Advertisement</span>
							<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<!-- 300x250 -->
<ins class="adsbygoogle"
     style="display:inline-block;width:300px;height:250px"
     data-ad-client="ca-pub-6883188387034598"
     data-ad-slot="4286918273"></ins>
<script>
(adsbygoogle = window.adsbygoogle || []).push({});
</script>						</div><!--mvp-flex-ad-->
					</div><!--mvp-flex-side-wrap-->
				</div><!--mvp-flex-side-out-->
					</div><!--mvp-widget-flex-wrap-->

		</div></section>			</div><!--mvp-home-widget-wrap-->
			</div><!--mvp-main-body-wrap-->
			<footer id="mvp-foot-wrap" class="left relative">
				<div id="mvp-foot-top" class="left relative">
					<div class="mvp-main-box">
						<div id="mvp-foot-logo" class="left relative">
															<a href="http://cronio.sv/"><img src="http://cronio.sv/wp-content/uploads/2018/03/logo-portada-3.png" alt="Diario Digital Cronio de El Salvador" data-rjs="2" /></a>
													</div><!--mvp-foot-logo-->
						<div id="mvp-foot-soc" class="left relative">
							<ul class="mvp-foot-soc-list left relative">
																	<li><a href="https://www.facebook.com/croniosv/" target="_blank" class="fa fa-facebook fa-2"></a></li>
																									<li><a href="https://twitter.com/croniosv" target="_blank" class="fa fa-twitter fa-2"></a></li>
																																	<li><a href="https://www.instagram.com/croniosv/" target="_blank" class="fa fa-instagram fa-2"></a></li>
																																	<li><a href="https://www.youtube.com/channel/UC9uaphREcIxCZHQgmoxkn0g/videos?disable_polymer=1" target="_blank" class="fa fa-youtube-play fa-2"></a></li>
																															</ul>
						</div><!--mvp-foot-soc-->
						<div id="mvp-foot-menu-wrap" class="left relative">
							<div id="mvp-foot-menu" class="left relative">
															</div><!--mvp-foot-menu-->
						</div><!--mvp-foot-menu-wrap-->
					</div><!--mvp-main-box-->
				</div><!--mvp-foot-top-->
				<div id="mvp-foot-bot" class="left relative">
					<div class="mvp-main-box">
						<div id="mvp-foot-copy" class="left relative">
							<p>Copyright © 2018 Diario Digital Cronio</p>
						</div><!--mvp-foot-copy-->
					</div><!--mvp-main-box-->
				</div><!--mvp-foot-bot-->
			</footer>
		</div><!--mvp-site-main-->
	</div><!--mvp-site-wall-->
</div><!--mvp-site-->
<div class="mvp-fly-top back-to-top">
	<i class="fa fa-angle-up fa-3"></i>
</div><!--mvp-fly-top-->
<div class="mvp-fly-fade mvp-fly-but-click">
</div><!--mvp-fly-fade-->
<script type="text/javascript">/* <![CDATA[ */ jQuery(document).ready( function() { jQuery.post( "http://cronio.sv/wp-admin/admin-ajax.php", { action : "entry_views", _ajax_nonce : "b905d38860", post_id : 17 } ); } ); /* ]]> */</script>
<link rel='stylesheet' id='svc-port-block-css-css'  href='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-block/css/css.css?ver=4.9.4' type='text/css' media='all' />
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-team/../assets/js/bootstrap.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-team/../assets/js/bootstrap-hover-dropdown.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/js/imagesloaded.pkgd.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-woo/../assets/js/owl.carousel.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/wp-all-in-one-grid/inc-team/../assets/js/custom.js?ver=4.9.4'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var impression_object = {"ajax_url":"http:\/\/cronio.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/adrotate/library/jquery.adrotate.dyngroup.js'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var click_object = {"ajax_url":"http:\/\/cronio.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type='text/javascript' src='http://cronio.sv/wp-content/plugins/adrotate/library/jquery.adrotate.clicktracker.js'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/themes/zox-news/js/mvpcustom.js?ver=4.9.4'></script>
<script type='text/javascript'>
	jQuery(document).ready(function($) {
	$(window).load(function(){
	var leaderHeight = $("#mvp-leader-wrap").outerHeight();
	var logoHeight = $("#mvp-main-nav-top").outerHeight();
	var botHeight = $("#mvp-main-nav-bot").outerHeight();
	var navHeight = $("#mvp-main-head-wrap").outerHeight();
	var headerHeight = navHeight + leaderHeight;
	var aboveNav = leaderHeight + logoHeight;
	var totalHeight = logoHeight + botHeight;
	var previousScroll = 0;
	$(window).scroll(function(event){
			var scroll = $(this).scrollTop();
			if ($(window).scrollTop() > aboveNav){
				$("#mvp-main-nav-top").addClass("mvp-nav-small");
				$("#mvp-main-nav-bot").css("margin-top", logoHeight );
			} else {
				$("#mvp-main-nav-top").removeClass("mvp-nav-small");
				$("#mvp-main-nav-bot").css("margin-top","0");
			}
			if ($(window).scrollTop() > headerHeight){
				$("#mvp-main-nav-top").addClass("mvp-fixed");
				$("#mvp-main-nav-bot").addClass("mvp-fixed1");
				$("#mvp-main-body-wrap").css("margin-top", totalHeight );
				$("#mvp-main-nav-top").addClass("mvp-fixed-shadow");
				$(".mvp-fly-top").addClass("mvp-to-top");
	    		if(scroll < previousScroll) {
					$("#mvp-main-nav-bot").addClass("mvp-fixed2");
					$("#mvp-main-nav-top").removeClass("mvp-fixed-shadow");
				} else {
					$("#mvp-main-nav-bot").removeClass("mvp-fixed2");
					$("#mvp-main-nav-top").addClass("mvp-fixed-shadow");
				}
			} else {
				$("#mvp-main-nav-top").removeClass("mvp-fixed");
				$("#mvp-main-nav-bot").removeClass("mvp-fixed1");
				$("#mvp-main-nav-bot").removeClass("mvp-fixed2");
				$("#mvp-main-body-wrap").css("margin-top","0");
				$("#mvp-main-nav-top").removeClass("mvp-fixed-shadow");
	    		$(".mvp-fly-top").removeClass("mvp-to-top");
			}
			previousScroll = scroll;
	});
	});
	});
	

	jQuery(document).ready(function($) {
	// Mobile Social Buttons More
	$(window).load(function(){
 		$(".mvp-soc-mob-right").on("click", function(){
			$("#mvp-soc-mob-wrap").toggleClass("mvp-soc-mob-more");
  		});
  	});
	});
  	

	jQuery(document).ready(function($) {
	$(window).load(function(){
		var leaderHeight = $("#mvp-leader-wrap").outerHeight();
		$("#mvp-site-main").css("margin-top", leaderHeight );
  	});

	$(window).resize(function(){
		var leaderHeight = $("#mvp-leader-wrap").outerHeight();
		$("#mvp-site-main").css("margin-top", leaderHeight );
	});

	});
  	

	jQuery(document).ready(function($) {
	$(".menu-item-has-children a").click(function(event){
	  event.stopPropagation();
	  location.href = this.href;
  	});

	$(".menu-item-has-children").click(function(){
    	  $(this).addClass("toggled");
    	  if($(".menu-item-has-children").hasClass("toggled"))
    	  {
    	  $(this).children("ul").toggle();
	  $(".mvp-fly-nav-menu").getNiceScroll().resize();
	  }
	  $(this).toggleClass("tog-minus");
    	  return false;
  	});

	// Main Menu Scroll
	$(window).load(function(){
	  $(".mvp-fly-nav-menu").niceScroll({cursorcolor:"#888",cursorwidth: 7,cursorborder: 0,zindex:999999});
	});
	});
	

	jQuery(document).ready(function($) {
	$(".infinite-content").infinitescroll({
	  navSelector: ".mvp-nav-links",
	  nextSelector: ".mvp-nav-links a:first",
	  itemSelector: ".infinite-post",
	  errorCallback: function(){ $(".mvp-inf-more-but").css("display", "none") }
	});
	$(window).unbind(".infscr");
	$(".mvp-inf-more-but").click(function(){
   		$(".infinite-content").infinitescroll("retrieve");
        	return false;
	});
	$(window).load(function(){
		if ($(".mvp-nav-links a").length) {
			$(".mvp-inf-more-but").css("display","inline-block");
		} else {
			$(".mvp-inf-more-but").css("display","none");
		}
	});
	});
	
</script>
<script type='text/javascript' src='http://cronio.sv/wp-content/themes/zox-news/js/scripts.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/themes/zox-news/js/retina.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-content/themes/zox-news/js/jquery.infinitescroll.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-includes/js/comment-reply.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://cronio.sv/wp-includes/js/wp-embed.min.js?ver=4.9.4'></script>
<!-- AdRotate JS -->
<script type="text/javascript">
jQuery(document).ready(function(){
if(jQuery.fn.gslider) {
	jQuery('.g-1').gslider({ groupid: 1, speed: 6000 });
}
});
</script>
<!-- /AdRotate JS -->

</body>
</html>