<!DOCTYPE html>
<html lang="en" dir="ltr" prefix="content: http://purl.org/rss/1.0/modules/content/  dc: http://purl.org/dc/terms/  foaf: http://xmlns.com/foaf/0.1/  og: http://ogp.me/ns#  rdfs: http://www.w3.org/2000/01/rdf-schema#  schema: http://schema.org/  sioc: http://rdfs.org/sioc/ns#  sioct: http://rdfs.org/sioc/types#  skos: http://www.w3.org/2004/02/skos/core#  xsd: http://www.w3.org/2001/XMLSchema# ">
  <head>
    <meta charset="utf-8" />
<script>(function(i,s,o,g,r,a,m){i["GoogleAnalyticsObject"]=r;i[r]=i[r]||function(){(i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)})(window,document,"script","https://www.google-analytics.com/analytics.js","ga");ga("create", "UA-19755360-7", {"cookieDomain":"auto"});ga("set", "anonymizeIp", true);ga("send", "pageview");</script>
<meta name="Generator" content="Drupal 8 (https://www.drupal.org)" />
<meta name="MobileOptimized" content="width" />
<meta name="HandheldFriendly" content="true" />
<meta name="viewport" content="width=device-width, initial-scale=1.0" />
<link rel="shortcut icon" href="/themes/custom/asam/favicon.ico" type="image/vnd.microsoft.icon" />
<script>window.a2a_config=window.a2a_config||{};a2a_config.callbacks=a2a_config.callbacks||[];a2a_config.templates=a2a_config.templates||{};a2a_config.no_3p=1;</script>

    <title>Home | Asamblea Legislativa de El Salvador</title>
    <style media="all">
@import url("/core/assets/vendor/normalize-css/normalize.css?p5legk");
@import url("/core/themes/stable/css/system/components/ajax-progress.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/align.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/autocomplete-loading.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/fieldgroup.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/container-inline.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/clearfix.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/details.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/hidden.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/item-list.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/js.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/nowrap.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/position-container.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/progress.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/reset-appearance.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/resize.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/sticky-header.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/system-status-counter.css?p5legk");
@import url("/core/themes/stable/css/system/components/system-status-report-counters.css?p5legk");
@import url("/core/themes/stable/css/system/components/system-status-report-general-info.css?p5legk");
@import url("/core/themes/stable/css/system/components/tabledrag.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/tablesort.module.css?p5legk");
@import url("/core/themes/stable/css/system/components/tree-child.module.css?p5legk");
@import url("/libraries/fontawesome/css/font-awesome.min.css?p5legk");
@import url("/core/themes/stable/css/views/views.module.css?p5legk");
@import url("/modules/addtoany/css/addtoany.css?p5legk");
@import url("/modules/asamblea_contenidos/css/asamblea-shortcodes.css?p5legk");
@import url("/modules/asamblea_social_media/css/asamblea-social-media.css?p5legk");
@import url("/modules/asamblea_social_media/soundmanager/css/bar-ui.css?p5legk");
@import url("/modules/asamblea_social_media/flowplayer-old/recursos/css.css?p5legk");
@import url("/libraries/bootstrap/css/bootstrap.css?p5legk");
</style>
<style media="all">
@import url("/core/themes/classy/css/components/action-links.css?p5legk");
@import url("/core/themes/classy/css/components/breadcrumb.css?p5legk");
@import url("/core/themes/classy/css/components/button.css?p5legk");
@import url("/core/themes/classy/css/components/collapse-processed.css?p5legk");
@import url("/core/themes/classy/css/components/container-inline.css?p5legk");
@import url("/core/themes/classy/css/components/details.css?p5legk");
@import url("/core/themes/classy/css/components/exposed-filters.css?p5legk");
@import url("/core/themes/classy/css/components/field.css?p5legk");
@import url("/core/themes/classy/css/components/form.css?p5legk");
@import url("/core/themes/classy/css/components/icons.css?p5legk");
@import url("/core/themes/classy/css/components/inline-form.css?p5legk");
@import url("/core/themes/classy/css/components/item-list.css?p5legk");
@import url("/core/themes/classy/css/components/link.css?p5legk");
@import url("/core/themes/classy/css/components/links.css?p5legk");
@import url("/core/themes/classy/css/components/menu.css?p5legk");
@import url("/core/themes/classy/css/components/more-link.css?p5legk");
@import url("/core/themes/classy/css/components/pager.css?p5legk");
@import url("/core/themes/classy/css/components/tabledrag.css?p5legk");
@import url("/core/themes/classy/css/components/tableselect.css?p5legk");
@import url("/core/themes/classy/css/components/tablesort.css?p5legk");
@import url("/core/themes/classy/css/components/tabs.css?p5legk");
@import url("/core/themes/classy/css/components/textarea.css?p5legk");
@import url("/core/themes/classy/css/components/ui-dialog.css?p5legk");
@import url("/core/themes/classy/css/components/messages.css?p5legk");
@import url("/themes/custom/asam/css/components/diputados.css?p5legk");
@import url("/themes/custom/asam/css/components/leyes-redes.css?p5legk");
@import url("/themes/custom/asam/css/components/node.css?p5legk");
@import url("/themes/custom/asam/css/components/identificadores.css?p5legk");
@import url("/themes/custom/asam/css/components/etiquetas.css?p5legk");
@import url("/themes/custom/asam/css/components/breadcrumb?p5legk");
@import url("/themes/custom/asam/css/components/menu.css?p5legk");
</style>
<style media="all">
@import url("/themes/custom/asam/css/components/style.css?p5legk");
@import url("/themes/custom/asam/css/components/dataTables.bootstrap.min.css?p5legk");
</style>

    
<!--[if lte IE 8]>
<script src="/core/assets/vendor/html5shiv/html5shiv.min.js?v=3.7.3"></script>
<![endif]-->

  </head>
  <body class="fontyourface path-frontpage">
        <a href="#main-content" class="visually-hidden focusable skip-link">
      Skip to main content
    </a>
    
        <section id="menuTop" class="makeMeSticky">
    <div  class="region region-top-header">
    <div id="block-asamblearedessocialesymediastreaming" class="block block-asamblea-social-media block-asamblea-social-media-block">
  
    
      
  <div id="menuTopContenedor">
    <div id="top-left-info" class="alignLeft">
      <div class="topBtnInicio"><a href="/"><img src="/modules/asamblea_social_media/images/icoAsamBlanco.svg" alt="Inicio"></a></div>
      <div class="topBtnTV">
        <a href="/asamblea-social-media/tv-player-popup" onclick="javascript:void window.open('/asamblea-social-media/tv-player-popup','1511189788195','width=800,height=600,toolbar=0,menubar=0,location=0,status=0,scrollbars=0,resizable=0,left=0,top=0');return false;">
          <img src="/modules/asamblea_social_media/images/9tvl-ico.svg" alt="Televisión Legislativa">
        </a>
      </div>
      <div id="top-right-info" class="topBtnRadio">
        <a href="/asamblea-social-media/radio-player-popup" onclick="javascript:void window.open('/asamblea-social-media/radio-player-popup','1511189788195','width=300,height=250,toolbar=0,menubar=0,location=0,status=0,scrollbars=0,resizable=0,left=0,top=0');return false;">
          <img src="/modules/asamblea_social_media/images/rl-ico.svg" alt="Radio Legislativa">
        </a>
      </div>
    </div>
    <div class="alignRight">
      <section id="buscarTop">
         <i class="fa fa-search search-icon search-block-no-buttom" aria-hidden="true" id="asam-global-search"></i>
      </section>
      <section id="redes-sociales">
        <ul class="rs-content">          
                  <div class="vacio">Este campo no tiene parámetros</div>
                
                  <li><a href="http://www.facebook.com/asamblea.legislativa" target="_blank" class="facebook-icono"><i class="fa fa-facebook-square" aria-hidden="true"></i></a></li>
                
                  <li><a href="https://twitter.com/AsambleaSV" target="_blank" class="twitter-icono"><i class="fa fa-twitter-square" aria-hidden="true"></i></a></li>
        
                  <li><a href="http://www.youtube.com/user/asambleaelsalvador" target="_blank" class="youtube-icono"><i class="fa fa-youtube" aria-hidden="true"></i></a></li>
                
                  <li><a href="http://flikr.com/photos/asamblealegislativa" target="_blank" class="flickr-icono"><i class="fa fa-flickr" aria-hidden="true"></i></a></li>
                </ul>
      </section>
      <section id="transparencia">
        <a href="https://transparencia.asamblea.gob.sv/" target="_blank" class="transparencia">PORTAL DE TRANSPARENCIA</a>
      </section>    
    </div>
  </div>
  </div>

  </div>

</section>

<div class="layout-container background-container">

  <header role="banner">
    
    <div class="logoNavMenu">
      <section id="header">
          <div  class="region region-header">
    <div id="block-asam-branding" class="block block-system block-system-branding-block">
  
    
        <a href="/" title="Home" rel="home" class="site-logo">
      <img class="headerimg logo" src="/themes/custom/asam/logo.svg" alt="Home" />
    </a>
      </div>

  </div>

      </section>
            <section id="menuPrincipal">  <div  class="region region-primary-menu">
    <nav role="navigation" aria-labelledby="block-asam-main-menu-menu" id="block-asam-main-menu" class="block block-menu navigation menu--main">
            
        
      
					<nav class="navbar navbar-custom">
				<div class="container-fluid">
					<div class="navbar-header">
					  <button type="button" class="navbar-toggle collapsed" data-toggle="collapse" data-target="#asamblea-nav-main-menu-bar" aria-expanded="false">
						<span class="sr-only">Toggle navigation</span>
						<span class="icon-bar"></span>
						<span class="icon-bar"></span>
						<span class="icon-bar"></span>
					  </button>
					</div>

					<div class="collapse navbar-collapse" id="asamblea-nav-main-menu-bar">
					
						<ul class="nav navbar-nav">
																																			<li class="dropdown">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Asamblea&nbsp;
																			
										<span class="caret"></span>
																				</a>
																				<ul class="dropdown-menu multi-level">
																					      
																										<li>
										<a href="/asamblea/diputadas-y-diputados">Diputadas y Diputados</a>
									</li>
																																<li>
										<a href="/diputados">Pleno Legislativo</a>
									</li>
																																<li>
										<a href="/junta-directiva">Junta Directiva</a>
									</li>
																																									<li class="dropdown-submenu">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Representación&nbsp;
																				</a>
																				<ul class="dropdown-menu">
																					      
																										<li>
										<a href="/diputados-departamento">Por Departamento</a>
									</li>
																																<li>
										<a href="/grupos-parlamentarios">Por Grupo Parlamantario</a>
									</li>
																	  
										</ul>
									</li>
																																<li>
										<a href="/asamblea/historia">Historia</a>
									</li>
																																<li>
										<a href="/asamblea/reglamento-interior">Reglamento Interior</a>
									</li>
																	  
										</ul>
									</li>
																																									<li class="dropdown">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Legislación&nbsp;
																			
										<span class="caret"></span>
																				</a>
																				<ul class="dropdown-menu multi-level">
																					      
																										<li>
										<a href="/legislacion/constitucion">Constitución</a>
									</li>
																																<li>
										<a href="/legislacion/anuarios-legislativos">Anuarios Legislativos</a>
									</li>
																																<li>
										<a href="/decretos/aniosdecretos">Decretos por Año</a>
									</li>
																																<li>
										<a href="/decretos/materiasgenero">Igualdad de Género</a>
									</li>
																	  
										</ul>
									</li>
																																									<li class="dropdown">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Sesión Plenaria&nbsp;
																			
										<span class="caret"></span>
																				</a>
																				<ul class="dropdown-menu multi-level">
																					      
																										<li>
										<a href="/agenda-legislativa/agenda">Agenda de Sesión Plenaria</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/asistencia-plenaria">Lista de Asistencia</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/notificaciones">Notificaciones</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/informes-trimestral">Informes de Comisiones</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/dictamenes">Dictámenes</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/correspondencia">Correspondencia</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/votaciones">Votaciones</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/convocatorias">Convocatoria</a>
									</li>
																																<li>
										<a href="/agenda-legislativa/resumen-plenaria">Resumen de la Sesión Plenaria</a>
									</li>
																																<li>
										<a href="/sesion-plenaria/archivo-historico">Archivo Histórico</a>
									</li>
																	  
										</ul>
									</li>
																																									<li class="dropdown">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Prensa&nbsp;
																			
										<span class="caret"></span>
																				</a>
																				<ul class="dropdown-menu multi-level">
																					      
																										<li>
										<a href="/asamblea-social-media/tv-player">TV Legislativa</a>
									</li>
																																<li>
										<a href="/asamblea-social-media/radio-player">Radio Legislativa</a>
									</li>
																																<li>
										<a href="/prensa/noticias">Últimas Noticias</a>
									</li>
																	  
										</ul>
									</li>
																																									<li class="dropdown">
																			<a href="" class="dropdown-toggle" data-toggle="dropdown" role="button" aria-haspopup="true" aria-expanded="false">Participación&nbsp;
																			
										<span class="caret"></span>
																				</a>
																				<ul class="dropdown-menu multi-level">
																					      
																										<li>
										<a href="/contact/consulta_ciudadana">Consulta Ciudadana</a>
									</li>
																																<li>
										<a href="/directorio-diputados">Directorio Parlamentario</a>
									</li>
																																<li>
										<a href="/participacion/oficinas-departamentales">Oficinas Departamentales</a>
									</li>
																	  
										</ul>
									</li>
																							</ul>
					</div>
				</div>
			</nav>
		  


  </nav>

  </div>
</section>
    </div>
  </header>
  <main role="main" class="main">
    
    <a id="main-content" tabindex="-1"></a>    
      <div  class="region region-carousel">
    <div class="block">
  
  
      <div id="diba-carousel" class="carousel slide" data-ride="carousel">
      <ol class="carousel-indicators">
                      <li data-target="#diba-carousel" data-slide-to="0" class = "active"></li>
                      <li data-target="#diba-carousel" data-slide-to="1" ></li>
                      <li data-target="#diba-carousel" data-slide-to="2" ></li>
                      <li data-target="#diba-carousel" data-slide-to="3" ></li>
                      <li data-target="#diba-carousel" data-slide-to="4" ></li>
            </ol>
      <ul class="carousel-inner" role="listbox">
                            <li class = "item active">
                          <img src="/sites/default/files/2018-03/NOTA%20HACIENDA-%20FOTO%20TITO.JPG" alt="  60 días de prórroga  para regular situación tributaria sin cobro de intereses " width="4155" height="2276">
                        <div class="carousel-caption">
                              <h2 class="caption-title">
                                      <a href="/node/6852">  60 días de prórroga  para regular situación tributaria sin cobro de intereses </a>
                                  </h2>
                                        </div>
          </li>
                            <li class = "item">
                          <img src="/sites/default/files/2018-03/NOTA%202-%20FOT%20GABY.JPG" alt="Aseguran fondos para pago de bonificación a los agentes de seguridad " width="3994" height="1796">
                        <div class="carousel-caption">
                              <h2 class="caption-title">
                                      <a href="/node/6854">Aseguran fondos para pago de bonificación a los agentes de seguridad </a>
                                  </h2>
                                        </div>
          </li>
                            <li class = "item">
                          <img src="/sites/default/files/2018-03/5E2A0296.JPG" alt="Presidente Guillermo Gallegos se reúne con el presidente de la Cámara de Representantes de Puerto Rico  " width="4998" height="3402">
                        <div class="carousel-caption">
                              <h2 class="caption-title">
                                      <a href="/node/6851">Presidente Guillermo Gallegos se reúne con el presidente de la Cámara de Representantes de Puerto Rico  </a>
                                  </h2>
                                        </div>
          </li>
                            <li class = "item">
                          <img src="/sites/default/files/2018-03/5E2A0535.JPG" alt="Asamblea Legislativa  otorga distinción honorífica “ Noble Amiga de El Salvador” a la embajadora de Chile " width="4317" height="3572">
                        <div class="carousel-caption">
                              <h2 class="caption-title">
                                      <a href="/node/6853">Asamblea Legislativa  otorga distinción honorífica “ Noble Amiga de El Salvador” a la embajadora de Chile </a>
                                  </h2>
                                        </div>
          </li>
                            <li class = "item">
                          <img src="/sites/default/files/2018-03/nota%20san%20vicente.jpg" alt="Asamblea Legislativa y Cruz Roja organizan taller sobre Primeros Auxilios en San Miguel" width="2000" height="800">
                        <div class="carousel-caption">
                              <h2 class="caption-title">
                                      <a href="/node/6850">Asamblea Legislativa y Cruz Roja organizan taller sobre Primeros Auxilios en San Miguel</a>
                                  </h2>
                                        </div>
          </li>
              </ul>
    <!-- Controls -->
    <a class="left carousel-control" href="#diba-carousel" role="button" data-slide="prev">
      <span class="glyphicon glyphicon-chevron-left" aria-hidden="true"></span>
      <span class="sr-only">Previous</span>
    </a>
    <a class="right carousel-control" href="#diba-carousel" role="button" data-slide="next">
      <span class="glyphicon glyphicon-chevron-right" aria-hidden="true"></span>
      <span class="sr-only">Next</span>
    </a>
    </div>
    

  
</div>

  </div>

      <div  class="region region-accesos-recursos">
    <div id="block-asambleaaccesosyrecursosblock" class="block block-asamblea-contenidos block-asamblea-accesos-recursos-block">
  
    
      <section class="accessSectionMain">
	<section class="row">
                            <!-- <div class="accessBox enlaces-x4"> -->
                <div class="accessBox col-lg-3 col-md-3 col-sm-6 col-xs-12">
                    <a class="accesBoxLinkContent" href="/leyes-decretos">
                        <h2>Leyes &raquo;</h2>
                    </a>
                    <div>
                        Búsqueda rápida de leyes, decretos o acuerdos, publicados en el Diario Oficial. Conoce también el proceso de Formación de Ley.
                    </div>
                </div>
                            <!-- <div class="accessBox enlaces-x4"> -->
                <div class="accessBox col-lg-3 col-md-3 col-sm-6 col-xs-12">
                    <a class="accesBoxLinkContent" href="/comisiones-legislativas">
                        <h2>Comisiones &raquo;</h2>
                    </a>
                    <div>
                        Conformados por Diputadas y Diputados propietarios, con el propósito de estudiar, analizar y aprobar, o rechazar las diferentes iniciativas de ley que se presentan a la Asamblea Legislativa.
                    </div>
                </div>
                            <!-- <div class="accessBox enlaces-x4"> -->
                <div class="accessBox col-lg-3 col-md-3 col-sm-6 col-xs-12">
                    <a class="accesBoxLinkContent" href="/prensa/noticias">
                        <h2>Noticias &raquo;</h2>
                    </a>
                    <div>
                        Noticias relacionadas con todo el que hacer parlamentario y toda la actividad en las diferentes comisiones legislativas.
                    </div>
                </div>
                            <!-- <div class="accessBox enlaces-x4"> -->
                <div class="accessBox col-lg-3 col-md-3 col-sm-6 col-xs-12">
                    <a class="accesBoxLinkContent" href="/enlaces">
                        <h2>Enlaces / Recursos &raquo;</h2>
                    </a>
                    <div>
                        Enlaces a diferentes recursos e información relacionados con la Asamblea Legislativa.
                    </div>
                </div>
            	</section>
    
</section>

  </div>

  </div>

      <div  class="region region-leyes-redes">
    <div id="block-asambleaultimosdecretos" class="block block-comisiones block-comisiones-ultimos-decretos-block">
  
    
      <div class="row-fluid">
                    <div class="col-lg-8 col-md-8 col-sm-6 col-xs-12 no-padding-left no-padding-right">
                                <div class="row-fluid">
                    <div class="col-sm-8 no-padding-left no-padding-right">
                                        <section>
    <div class="tituloLeyesFront">Últimos decretos</div>
    <div class="leyesFrontBox">
        <div class="panel panel-default">
            <div class="panel-body">
                <ul class="News leyesFrontList">
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3371">
                                924&nbsp;-&nbsp;EXONÉRASE DEL PAGO DE IMPUESTOS, A LEAGUE C.A., LIMITADA DE C.V. DE LA DONACIÓN DE UN COMPRESOR DE AIRE, Y UN SECADOR DE AIRE REFRIGERADO, A FAVOR DE LA DIRECCIÓN GENERAL DE CENTROS PENALES.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3372">
                                925&nbsp;-&nbsp;PRORROGASE LA LEY TRANSITORIA PARA FACILITAR EL CUMPLIMIENTO VOLUNTARIO DE OBLIGACIONES TRIBUTARIAS Y ADUANERAS.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3335">
                                921&nbsp;-&nbsp;Refórmase la Ley de Presupuesto, en la parte correspondiente a los Ramos de Relaciones Exteriores, Fiscalía General de la República y Registro Nacional de las Personas Naturales (para el Tribunal Supremo Electoral), para incorporar $3,289,000.00.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3352">
                                913&nbsp;-&nbsp;LEY DE CREACIÓN DEL INSTITUTO NACIONAL DE FORMACIÓN DOCENTE.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3353">
                                914&nbsp;-&nbsp;LEY ESPECIAL REGULADORA PARA LA CONTRATACIÓN Y COLOCACIÓN DE LA GENTE DE MAR EN BUQUES DE BANDERA EXTRANJERA.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3354">
                                915&nbsp;-&nbsp;AUTORÍZASE EL INGRESO, TRÁNSITO Y ESTACIONAMIENTO EN AGUAS TERRITORIALES, DE LA FLOTA DE LA FUERZA NAVAL DE LA REPÚBLICA DE CHINA (TAIWÁN).
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3355">
                                916&nbsp;-&nbsp;REFORMA A LA LEY DE CONTROL Y REGULACIÓN DE ARMAS, MUNICIONES, EXPLOSIVOS Y ARTÍCULOS SIMILARES.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3357">
                                917&nbsp;-&nbsp;REFÓRMASE LA LEY DE PRESUPUESTO, EN LA PARTE QUE CORRESPONDE AL RAMO DE EDUCACIÓN, PARA INCORPORAR $6,257,154.00.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3358">
                                918&nbsp;-&nbsp;REFÓRMASE LA LEY DE SALARIOS EN LA PARTE CORRESPONDIENTE AL ESCALAFÓN DE LA UNIVERSIDAD DE EL SALVADOR; PARA BENEFICIAR A 3,493 PLAZAS DE LEY DE SALARIOS.
                            </a>
                        </li>
                                            <li class="news-item">
                            <a href="https://www.asamblea.gob.sv//decretos/details/3360">
                                919&nbsp;-&nbsp;REFÓRMASE EL D.L. 880/2018.
                            </a>
                        </li>
                                    </ul>
            </div>
            <div class="panel-footer"> </div>
        </div>
    </div>
</section>
<input type="hidden" id="asamblea_ultimos_decretos_cantidad" value="10">
                                   </div>
                   <div class="col-sm-4 no-padding-left no-padding-right">
                        <section>
                            <div class="tituloBusquedaFront">Búsqueda de leyes</div>
                            <div class="busquedaFrontBox">
                                <form class="form-horizontal col-md-12" id="block-mini-busqueda-form" action="https://www.asamblea.gob.sv/decretos/resultadobusqueda/" method="get">
        <div class="input-group" id="block-mini-busqueda-palabra-interes-wrapper">
            <span class="input-group-addon">
                <span class="glyphicon glyphicon-search col-md-1" aria-hidden="true"></span>
            </span>
            <input type="text" class="form-control input-sm" id="block-mini-busqueda-palabra-interes" placeholder="Búsqueda de Leyes y Decrétos" name="palabras_interes" />
        </div>
        <div id="block-mini-busqueda-tipo-documento">
            <div><input type="checkbox" name="tiposdecreto[]" value="2C7F9863-ACD6-4D66-B520-1A61DEC2A207"><span>Código</span></div>
            <div><input type="checkbox" name="tiposdecreto[]" value="93F5C05D-30B9-4779-84F6-67E61C1911CD"><span>Decreto</span></div>
            <div><input type="checkbox" name="tiposdecreto[]" checked="checked" value="597D1D4D-DA66-4878-A841-3D08AD6723F6"><span>Ley</span></div>
            <div><input type="checkbox" name="tiposdecreto[]" value="E892660B-B733-426D-BF2D-059D12CFFDCB"><span>Reglamento</span></div>
        </div>
        <input class="btn btn-default col-md-12" id="block-mini-busqueda-boton-buscar" type="submit" value="Buscar">
</form>
<p class="busqueda-texto-info">El contenido de este servicio se encuentra en permanente actualización por la Unidad de Índice Legislativo, por lo que de no encontrar el documento requerido lo puede solicitar a los teléfonos 2281-9225, 2281-9299 y 2281-9228 o al correo electrónico <a href="mailto:indice.legislativo@asamblea.gob.sv">indice.legislativo@asamblea.gob.sv</a>.</p>
<a class="btn btn-info col-md-12" id="block-mini-busqueda-link-busqueda-avanzada" href="https://www.asamblea.gob.sv/decretos/busquedadecretos">Búsqueda avanzada</a>   
                            </div>
                            
                        </section>
                   </div>
                </div>
                            </div>
            <div class="col-lg-4 col-md-4 col-sm-6 col-xs-12 no-padding-left no-padding-right">
                <section>
    <div class="tituloRedesFront">Nuestras redes</div>
    <div class="redesFrontBox">
        <ul class="nav nav-tabs" id="social-asamblea-tabs">
            <li class="active">
                <a data-toggle="tab" href="#twitter-asamblea">Últimos tweets</a>
            </li>
            <li>
                <a data-toggle="tab" href="#facebook-asamblea">Últimos post</a>
            </li>
        </ul>
        <div class="tab-content" id="social-asamblea-tabs-content">
            <div id="twitter-asamblea" class="tab-pane fade in active scrollRedes">
                <a class="twitter-timeline" data-lang="es" data-dnt="true" href="https://twitter.com/AsambleaSV?ref_src=twsrc%5Etfw">
                    
                </a>
                <script async src="//platform.twitter.com/widgets.js" charset="utf-8"></script>
            </div>
            <div id="facebook-asamblea" class="tab-pane fade scrollRedes">
                <iframe
                    id="iframe-facebook-asamblea"
                    src="https://www.facebook.com/plugins/page.php?href=https://www.facebook.com/asamblea.legislativa&tabs=timeline&width=450&height=345&small_header=true&adapt_container_width=true&hide_cover=true&show_facepile=false&appId"
                    width="100%"
                    height="346"
                    style="border:none;overflow:hidden"
                    scrolling="no"
                    frameborder="0"
                    allowTransparency="true">

                </iframe>
            </div>
        </div>
    </div>                
</section>
            </div>
        </div>
  </div>

  </div>

    <div class="layout-content">

      <div class="container-fluid">
        
        
        
        <section class="row-fluid">
                      <div class="col-md-12">
                  <div  class="region region-content">
    <div class="views-element-container"><div class="view view-duplicate-of-frontpage view-id-duplicate_of_frontpage view-display-id-page_1 js-view-dom-id-d9e510f864312f9ea4f8c335b6b61bcbe46f1368518bdc85a882f7335f167a83">
  
    
      
  
      
          </div>
</div>

  </div>

                <span class="a2a_kit a2a_kit_size_32 addtoany_list"></span>
            </div>
                  </section>        
      </div>

    </div>    
  </main>

      <footer role="contentinfo">
        <div  class="region region-footer">
    <div id="block-footerestatico" class="block block-block-content block-block-content6756111a-9201-4f14-8014-bfcf7f0221f1">
  
    
      
            <div class="clearfix text-formatted field field--name-body field--type-text-with-summary field--label-hidden field__item"><footer><!-- FONDO PARTICULAS --><!-- div id="particles-js">&nbsp;</div --><!-- FIN FONDO PARTICULAS --><div class="row-fluid footer-info">
<div class="col-lg-4 col-md-4 col-sm-4 col-xs-12 no-padding-left no-padding-right">
<h5>Oficina de Información Pública</h5>

<p><b>Teléfonos:</b><br />
(503) 2281 – 9382<br /><b>Correos Electrónico:</b><br /><a href="mailto:transparencia@asamblea.gob.sv">transparencia@asamblea.gob.sv</a></p>
</div>

<div class="col-lg-4 col-md-4 col-sm-4 col-xs-12 no-padding-left no-padding-right footer-logo"><img alt="footer" class="footerImg" src="https://www.asamblea.gob.sv/themes/custom/asam/images/footer.svg" /></div>

<div class="col-lg-4 col-md-4 col-sm-4 col-xs-12 no-padding-left no-padding-right">
<h5>Oficina de Índice Legislativo</h5>

<p><b>Teléfonos:</b><br />
(503) 2281 - 9225<br />
(503) 2281 - 9299<br />
(503) 2281 - 9228<br />
 <br />
 <br /><b>Correo electrónico:</b><br /><a href="mailto:indice.legislativo@asamblea.gob.sv">indice.legislativo@asamblea.gob.sv</a></p>
</div>
</div>

<div class="row-fluid">
<div class="col-md-12">
<p class="dirpostal">Centro de Gobierno "José Simeón Cañas", Palacio Legislativo, San Salvador, El Salvador. CP 1101 Teléfono: 2281-9000.</p>
</div>
</div>
</footer></div>
      
  </div>

  </div>

    </footer>
  
</div>
    <script type="application/json" data-drupal-selector="drupal-settings-json">{"path":{"baseUrl":"\/","scriptPath":null,"pathPrefix":"","currentPath":"node","currentPathIsAdmin":false,"isFront":true,"currentLanguage":"en"},"pluralDelimiter":"\u0003","google_analytics":{"trackOutbound":true,"trackMailto":true,"trackDownload":true,"trackDownloadExtensions":"7z|aac|arc|arj|asf|asx|avi|bin|csv|doc(x|m)?|dot(x|m)?|exe|flv|gif|gz|gzip|hqx|jar|jpe?g|js|mp(2|3|4|e?g)|mov(ie)?|msi|msp|pdf|phps|png|ppt(x|m)?|pot(x|m)?|pps(x|m)?|ppam|sld(x|m)?|thmx|qtm?|ra(m|r)?|sea|sit|tar|tgz|torrent|txt|wav|wma|wmv|wpd|xls(x|m|b)?|xlt(x|m)|xlam|xml|z|zip"},"user":{"uid":0,"permissionsHash":"24471894161de449c0e44e273731f6c9f72dea222ef16c27142a038cd2503832"}}</script>
<script src="/core/assets/vendor/domready/ready.min.js?v=1.0.8"></script>
<script src="/core/assets/vendor/jquery/jquery.min.js?v=3.2.1"></script>
<script src="/core/misc/drupalSettingsLoader.js?v=8.4.2"></script>
<script src="/core/misc/drupal.js?v=8.4.2"></script>
<script src="/core/misc/drupal.init.js?v=8.4.2"></script>
<script src="https://static.addtoany.com/menu/page.js" async></script>
<script src="/modules/addtoany/js/addtoany.js?v=8.4.2"></script>
<script src="/modules/asamblea_contenidos/js/asamblea-shortcodes.js?p5legk"></script>
<script src="/modules/asamblea_social_media/js/google-swfobject.js?p5legk"></script>
<script src="/modules/asamblea_social_media/js/asamblea-social-media.js?p5legk"></script>
<script src="/modules/asamblea_social_media/soundmanager/script/soundmanager2.js?p5legk"></script>
<script src="/modules/asamblea_social_media/soundmanager/script/bar-ui.js?p5legk"></script>
<script src="/modules/asamblea_social_media/flowplayer-old/recursos/flowplayer-3.2.6.min.js?p5legk"></script>
<script src="/modules/asamblea_social_media/flowplayer-old/recursos/9tvl.js?p5legk"></script>
<script src="/libraries/bootstrap/js/bootstrap.js?p5legk"></script>
<script src="/modules/google_analytics/js/google_analytics.js?v=8.4.2"></script>
<script src="/themes/custom/asam/js/bootstrap-search.js?v=2.x"></script>
<script src="/themes/custom/asam/js/add-img-responsive-class.js?v=2.x"></script>
<script src="/themes/custom/asam/js/dataTables.min.js?v=2.x"></script>
<script src="/themes/custom/asam/js/dataTables.bootstrap.min.js?v=2.x"></script>
<script src="/themes/custom/asam/js/jquery.touchSwipe.min.js?v=2.x"></script>
<script src="/themes/custom/asam/js/swipe.bootstrap.carousel.js?v=2.x"></script>
<script src="/themes/custom/asam/js/jquery.bootstrap.newsbox.js?v=2.x"></script>
<script src="/themes/custom/asam/js/news-home.newsbox.js?v=2.x"></script>

  </body>
</html>