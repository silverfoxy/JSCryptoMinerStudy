﻿<!DOCTYPE html>
<html lang="es" xmlns="http://www.w3.org/1999/xhtml">
<head>
	<meta charset="utf-8">
	<meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
	<meta name="viewport" content="width=device-width, initial-scale=1">
	<link rel="icon" type="image/x-icon" href="favicon.ico" />
	<title>Dirección de Educación Virtual de la Universidad Tecnológica de El Salvador</title>
	<meta name="Keywords" content="clases virtual, salon de apoyo, islas, el salvador, salvador, universidad, licenciatura, ingenieria, 
									asignatura, asignaturas, moodle, curso, ciclo  
									administracion virtual, carrera virtual, ingenieria virtual, mercadeo virtual, academico, profesor, unidades,
									edutec, educacion a distancia, utec, 
									universidad tecnologia, educacion a distancia el salvador, universidad tecnologica, EDUTEC, 
									semipresenciales, seminario taller utec, educacion a distancia utec" />
	<meta name="Description" content="EDUTEC - Educacion a Distancia de la Universidad Tecnologica de El Salvador, 
										A partir de junio del 2002 la Universidad Tecnolgica consolid el Proyecto de Educacin a Distancia, 
										creando el sitio EDUTEC, y generando con ello valiosos aportes al desarrollo nacional que amplan 
										el alcance de las comunidades acadmicas, y poniendo de manifiesto lo establecido en 
										la MISION y VISION de la Universidad Tecnologica de El Salvador." />
	<meta name="reply-to" content="utecvirtual@utec.edu.sv" />
	<meta name="title" content="Dirección de Educación Virtual de la Universidad Tecnológica de El Salvador"  />
	<meta name="author" content="UTECVIRTUAL"  />
	<meta name="Classification" content="Universidad" />
	<meta name="Language" content="Spanish, English, French, German, Italian, Chinese Simplified" />
	<meta name="copyright" content="UTECVIRTUAL" />
	<meta name="city" content="San Salvador" />
	<meta name="country" content="El Salvador" />
	<meta name="distribution" content="Global" />
	<meta name="Revisit-After" content="8 days" />

	<meta itemprop="name" content="Utec Virtual">
	<meta itemprop="description" content="Dirección de Educación Virtual de la Universidad Tecnológica de El Salvador">
	<meta itemprop="image" content="http://www.edutec.edu.sv/images/logo.png">

	<link rel="stylesheet" href="https://maxcdn.bootstrapcdn.com/font-awesome/4.5.0/css/font-awesome.min.css">
	<link rel='stylesheet' href='https://fonts.googleapis.com/css?family=Roboto:400,300,500'>
	<!-- Latest compiled and minified CSS -->
	<link rel="stylesheet" href="https://maxcdn.bootstrapcdn.com/bootstrap/3.3.6/css/bootstrap.min.css" integrity="sha384-1q8mTJOASx8j1Au+a5WDVnPi2lkFfwwEAa8hDDdjZlpLegxhjVME1fgjWPGmkzs7" crossorigin="anonymous">
	<!-- Cargaremos estilos moviles -->
	<link rel="stylesheet" media="only screen and (max-device-width: 480px) and (min-device-width: 320px)" href="css/mobile.css" type="text/css" />
	<link rel="stylesheet" media="handheld, only screen and (max-device-width: 319px)" href="css/mobile_simple.css" type="text/css" />
	<style>
	body {
		font-family: 'Roboto', sans-serif;
	}
	menuitem a {
		height:63px;
		display:inline-block;
		text-decoration:none;
		color:#000;
		padding:0 10px;
	}
	menuitem a:hover {
		background-color:#494949;
		color:#fff;
	}
	menuitem a.active {
		background-color:#494949;
		color:#fff;
	}
	div.float-form div.content-form
{
    background: #641A33;
    padding: 8px;
    padding-right: 0px;
    padding-bottom: 0px;
}

div.float-form-inner div.content-form
{
    background: #E8E8E8;
    padding: 8px;
    padding-right: 8px;
    padding-bottom: 0px;
    position: relative;
}

div.float-form-inner div.content-form input
{
    width: 240px;
    margin-bottom: 6px;
}

div.float-form-inner div.content-form select
{
    width: 254px;
    margin-bottom: 6px;
}

div.float-form-inner div.content-form a.close-equis
{
    position: absolute;
    right: -15px;
    top: -50px;
}
.no-padding {
	padding: 0;
}
.content-form {
	margin:0 auto;
	width:83%;
}
.content-form img {
	width: 100%;
}
/*
div.float-form
{
    left: 150px;
    position: absolute;
    top: 120px;
    width: 330px;
    z-index: 999;
}
*/
div.float-form-inner
{
    width: 270px;
    display: inline-block;
}
/*
.black_button {
	width: 90%;
    display: block;
    height: 60px;
    border: 0;
    background: #3c3c3c;
    color: white;
    font-size: 1.5em;
    text-align: left;
    line-height: 60px;
    padding-left: 1.5em;
    border-radius: 10px 10px 10px 10px;
    -moz-border-radius: 10px 10px 10px 10px;
    -webkit-border-radius: 10px 10px 10px 10px;
    border: 0px solid #000000;
    -webkit-box-shadow: 2px 4px 5px 1px rgba(0,0,0,0.75);
    -moz-box-shadow: 2px 4px 5px 1px rgba(0,0,0,0.75);
    box-shadow: 2px 4px 3px 1px rgba(0,0,0,0.75);
}
*/
.black_button {
    width: 90%;
    display: block;
    background: #3c3c3c;
    color: white;
    text-align: center;
    border-radius: 10px 10px 10px 10px;
    -moz-border-radius: 10px 10px 10px 10px;
    -webkit-border-radius: 25px;
    border: 0px solid #000000;
    -webkit-box-shadow: 2px 4px 5px 1px rgba(0,0,0,0.75);
    -moz-box-shadow: 2px 4px 5px 1px rgba(0,0,0,0.75);
    box-shadow: 2px 4px 3px 1px rgba(0,0,0,0.75);
    font-size: 1.1em;
    padding: 15px;
}

.black_button:hover {
	color: #a7a7a7;
    text-decoration: none;
    background: #4f4f4f;
}
.info_button {
	color: gainsboro;
    width: 85%;
    text-align: center;
    font-size: 0.9em;
    margin-bottom: 20px;
    padding-top: 6px;
}
.icon-space {
	width: 40px;
	height: 44px;
	float: left;
    margin-top: 10px;
    margin-right: 15px;
	background:url(img/sprite-home.png) -100px -500px #3c3c3c no-repeat;
}
.icon-info {
	background-position: 10px 0px;
}

.icon-req {
	background-position: -42px 0px;
}
.icon-hist {
	background-position: -92px 0px;
}
.icon-4x {
	font-size: 4em;
}
.icon-curso {
	background-position: -140px 0px;
}
   /* jssor slider bullet navigator skin 05 css */
        /*
        .jssorb05 div           (normal)
        .jssorb05 div:hover     (normal mouseover)
        .jssorb05 .av           (active)
        .jssorb05 .av:hover     (active mouseover)
        .jssorb05 .dn           (mousedown)
        */
        .jssorb05 {
            position: absolute;
        }
        .jssorb05 div, .jssorb05 div:hover, .jssorb05 .av {
            position: absolute;
            /* size of bullet elment */
            width: 16px;
            height: 16px;
            background: url('img/b05.png') no-repeat;
            overflow: hidden;
            cursor: pointer;
        }
        .jssorb05 div { background-position: -7px -7px; }
        .jssorb05 div:hover, .jssorb05 .av:hover { background-position: -37px -7px; }
        .jssorb05 .av { background-position: -67px -7px; }
        .jssorb05 .dn, .jssorb05 .dn:hover { background-position: -97px -7px; }

        .head-title {
        	font-size:2vw;
        }
		/* agregamos media query para texto footer */
		@media only screen and (max-width: 768px) {
			.head-title {
        		font-size:3vw;
        	}
        	.content-form {
				width:100%;
			}
		}
		@media only screen and (min-width: 1280px) {
        	.content-form {
				width:74%;
			}
			
		}
		@media only screen and (min-width: 1460px) {
        	.content-form {
				width:61%;
			}
			.content {
				max-height:370px;
			}
		}
		@media only screen and (max-width: 480px) {
			.content-form {
				width:100%;
			}
			.content {
				max-height:250px;
			}
			.content-form img {
				width: 100%;
			}
			.foot-form-solicitud {
				text-align:center;
			}
			.head-title {
        		font-size:5vw;
        	}
			  .col-ssx-1, .col-ssx-2, .col-ssx-3, .col-ssx-4, .col-ssx-5, .col-ssx-6, .col-ssx-7, .col-ssx-8, .col-ssx-9, .col-ssx-10, .col-ssx-11, .col-ssx-12 {
				float: left;
			  }
			  .col-ssx-12 {
				width: 100%;
			  }
			  .col-ssx-11 {
				width: 91.66666667%;
			  }
			  .col-ssx-10 {
				width: 83.33333333%;
			  }
			  .col-ssx-9 {
				width: 75%;
			  }
			  .col-ssx-8 {
				width: 66.66666667%;
			  }
			  .col-ssx-7 {
				width: 58.33333333%;
			  }
			  .col-ssx-6 {
				width: 50%;
			  }
			  .col-ssx-5 {
				width: 41.66666667%;
			  }
			  .col-ssx-4 {
				width: 33.33333333%;
			  }
			  .col-ssx-3 {
				width: 25%;
			  }
			  .col-ssx-2 {
				width: 16.66666667%;
			  }
			  .col-ssx-1 {
				width: 8.33333333%;
			  }
		}
		 .readmore + [data-readmore-toggle], .readmore[data-readmore]{display: block; margin: 15px;}
		 .readmore[data-readmore]{transition: height 75ms;overflow: hidden;}
		 .btns-v a {
		 	text-align: left;
		 	padding-left: 10px;
		 }
		 .btn-outline {
    background-color: transparent;
    color: inherit;
    transition: all .5s;
}

.btn-primary.btn-outline {
    color: #428bca;
}

.btn-success.btn-outline {
    color: #5cb85c;
}

.btn-info.btn-outline {
    color: #5bc0de;
}

.btn-warning.btn-outline {
    color: #f0ad4e;
}

.btn-danger.btn-outline {
    color: #d9534f;
}

.btn-primary.btn-outline:hover,
.btn-success.btn-outline:hover,
.btn-info.btn-outline:hover,
.btn-warning.btn-outline:hover,
.btn-danger.btn-outline:hover {
    color: #fff;
}
	</style>
	<link rel="stylesheet" href="css/sweetalert.css" type="text/css" />
	<!-- HTML5 shim and Respond.js for IE8 support of HTML5 elements and media queries -->
    <!--[if lt IE 9]>
      <script src="https://oss.maxcdn.com/html5shiv/3.7.2/html5shiv.min.js"></script>
      <script src="https://oss.maxcdn.com/respond/1.4.2/respond.min.js"></script>
    <![endif]-->
	<!-- Analytics -->
	<script>
	  (function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
	  (i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
	  m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
	  })(window,document,'script','//www.google-analytics.com/analytics.js','ga');
	  ga('create', 'UA-71894674-1', 'auto');
	  ga('send', 'pageview');
	</script>
</head>
<body>
	<!-- Google Tag Manager -->
	<noscript><iframe src="//www.googletagmanager.com/ns.html?id=GTM-W8JTJL"
	height="0" width="0" style="display:none;visibility:hidden"></iframe></noscript>
	<script>(function(w,d,s,l,i){w[l]=w[l]||[];w[l].push({'gtm.start':
	new Date().getTime(),event:'gtm.js'});var f=d.getElementsByTagName(s)[0],
	j=d.createElement(s),dl=l!='dataLayer'?'&l='+l:'';j.async=true;j.src=
	'//www.googletagmanager.com/gtm.js?id='+i+dl;f.parentNode.insertBefore(j,f);
	})(window,document,'script','dataLayer','GTM-W8JTJL');</script>
	<!-- End Google Tag Manager -->
	<!--[if lt IE 8]>
		<p class="chromeframe">Estas usando un navegador <strong>desactualizado</strong>. Por favor <a href="http://browsehappy.com/">Actualiza tu navegador</a> o <a href="http://www.google.com/chromeframe/?redirect=true">activa Google Chrome Frame</a> para mejorar la experiencia.</p>
	<![endif]-->
	<header style="background:url(images/header-bg.png) no-repeat;">
		<div id="logo" style="width:300px;padding:20px;margin-left:20px;">
			<img src="images/logo-utec.png" alt="Universidad Tecnologica de El Salvador" style="width:100%" />
		</div>
		 <nav class="navbar navbar-inverse" style="background:url(images/menu-bg.jpg) repeat-x; border:0;margin-bottom:0;">
		  <div class="container">
			<div class="navbar-header">
			  <button type="button" class="navbar-toggle collapsed" data-toggle="collapse" data-target="#navbar" aria-expanded="false" aria-controls="navbar">
				<span class="sr-only">Ver Enlaces</span>
				<span class="icon-bar"></span>
				<span class="icon-bar"></span>
				<span class="icon-bar"></span>
			  </button>
			  <a class="navbar-brand" href="/"><i class="fa fa-home fa-lg"></i></a>
			</div>
			<div id="navbar" class="collapse navbar-collapse">
			  <ul class="nav navbar-nav">
				<li><a target="_blank" href="http://www.utec.edu.sv/">UTEC</a></li>
				<li><a target="_blank" href="http://portal.utec.edu.sv/">PORTAL EDUCATIVO</a></li>
				<li><a target="_blank" href="http://www.utec.edu.sv/Inicio/Publicaciones">PUBLICACIONES</a></li>

					<script type="text/javascript" src="https://unpkg.com/sweetalert2@7.3.5/dist/sweetalert2.all.js"></script>
					<script src="bower_components/sweetalert2/dist/sweetalert2.min.js"></script>
					<link rel="stylesheet" href="bower_components/sweetalert2/dist/sweetalert2.min.css">
					<script type="text/javascript">
						function alerta() {
							swal({
		  						title: 'Nueva plataforma virtual',
		  						text: 'Para alumnos de la carrera virtual.',
		  						timer: 3000,
		  						type: 'info'
								});
						}
					</script>

				<style type="text/css">
				.coor_red{
							box-shadow: 0px 0px 15px #5d0a28;
							color: black !important;
						
						}
						.coor_red:hover{
							color: #5d0a28 !important;
							transition-property: color;
							transition-property: box-shadow;
							transition-duration: 0.9s !important;
							box-shadow: 0px 0px 35px #5d0a28;

						}

				</style>
				<li><a target="_blank" href="https://utds.mrooms.net/" class="coor_red"  onmouseleave="alerta()">CARRERAS VIRTUALES</a></li>
				<!-- <li><a href="http://lapalabra.utec.edu.sv/">LA PALABRA</a></li>
				<li><a href="http://www.graduadoutec.edu.sv/">INSTITUTO GRADUADOS</a></li>
				<li><a href="http://biblioteca.utec.edu.sv/">BIBLIOTECA UTEC</a></li> -->
			  </ul>
			</div><!--/.nav-collapse -->
		  </div>
		</nav>
		<div id="social" style="float:right;margin-right:30px;padding-right:8em;">
			<a href="https://plus.google.com/u/0/+UtecvirtualEduSv79" target="_blank" style="float:left;"><img src="../images/gp-social-icon.jpg" /></a>
			<a href="https://www.facebook.com/utecvirtual" target="_blank" style="float:left;"><img src="../images/fb-social-icon.jpg" /></a>
		</div>
		<div style="clear:both;"></div>
		<section id="login" style="background:url(images/login-bg.jpg) center center no-repeat; background-size:cover; width:100%;">
			<div id="jssor_1" style="position: relative; margin: 0 auto; top: 0px; left: 0px; width: 1300px; height: 313px; overflow: hidden; visibility: hidden;">
				<!-- Loading Screen -->
				<div data-u="loading" style="position: absolute; top: 0px; left: 0px;">
					<div style="filter: alpha(opacity=70); opacity: 0.7; position: absolute; display: block; top: 0px; left: 0px; width: 100%; height: 100%;"></div>
					<div style="position:absolute;display:block;background:url('img/loading.gif') no-repeat center center;top:0px;left:0px;width:100%;height:100%;"></div>
				</div>
				<div data-u="slides" style="cursor: default; position: relative; top: 0px; left: 0px; width: 1300px; height: 313px; overflow: hidden;">
					<div data-p="225.00" style="display: none;">
						<img data-u="image" src="img/portada01.jpg" alt="Portada 1" />
					</div>
					<div data-p="225.00" style="display: none;">
						<img data-u="image" src="img/portada02.jpg" alt="Portada 2" />
					</div>
					<div data-p="225.00" style="display: none;">
						<img data-u="image" src="img/portada03.jpg" alt="Portada 3" />
					</div>
					<div u='any' style='position: absolute; top: 10px; left: 795px; width: 100px; height: 26px;'>
						<div id="innerLogin" style="margin-right:20px;width:350px;">
							<div style="background:url(images/login.png) no-repeat;background-size:contain;padding:80px 20px; 40px">
							<form id="frmLogin" style="margin-top:5px;" name="frmLogin" action="acceso/login.php" method="post" onsubmit="return validar(this);">
								<input type="text" name="txtUser" id="txtUser" style="width:100%;height:40px;" maxlength="25" onkeydown="return alfanumerico(event,this);" placeholder="Usuario: Ej. 2200002016" />
								<br /><br />
								<input type="password" name="txtPass" id="txtPass" style="width:100%;height:40px;" maxlength="50" autocomplete="off" placeholder="Contrasena: Ej. **********" />
								<br /><br />
								<input type="submit" name="btnSubmit" id="btnSubmit" style="width:100%;height:50px;font-size:1.9em;color:#c9c9c9;background-color:#313131;border:0;" value="INGRESAR" />
							</form>
							</div>
						</div>
					</div>
				</div>
				<!-- Bullet Navigator -->
				<div data-u="navigator" class="jssorb05" style="bottom:16px;right:16px;" data-autocenter="1">
					<!-- bullet navigator item prototype -->
					<div data-u="prototype" style="width:16px;height:16px;"></div>
				</div>
			</div>
			
			<div style="clear:both;"></div>
		</section>
	</header>
	
	<section>
		<div class="container-fluid">
			<div class="row news-wrapper" style="width: 95%;margin: 5px auto;background-color: #e7e7e7;font-size: small;">
			  <div class="content" style="padding: 1% 5% 0.5%;">
				<div>
					<span style="font-weight: bold;color: #980A4D;">Noticias.</span>

			<!--<strong>Oportunidad de beca Estudiantes virtuales.</strong>La Dirección de Internacionalización Académica-DIA, &nbsp;de la Rectoría UNIMINUTO Virtual y a Distancia de la Corporación Universitaria Minuto de Dios –UNIMINUTO (Colombia), invita a las universidades internacionales aliadas, a participar de la convocatoria de becas de intercambio.-->


					<strong>A los alumnos de carreras no presenciales, les informamos que el ciclo 01-2018 cambiaremos de plataforma tecnológica, entérese ingresando a su área virtual.</strong>
				</div>
				<!-- <div style="text-align:right"><a href="./noticias.php?id=1001">Leer Mas →</a><a></a></div> -->
			  </div>
			</div>
			<div class="row">
				<div class="textHeader" style="font-size:1.5em; width:70%;margin:30px auto;text-align:center;color:#980A4D;">
					<h1 class="head-title">LA UNIVERSIDAD TECNOLÓGICA TE OFRECE CARRERAS VIRTUALES<br />PARA CONTINUAR CON TU PREPARACIÓN</h1>
				</div>
			</div>
			<div class="row">
				<div class="col-ssx-12 col-xs-6 col-sm-4">
					<div class="content readmore1">
						<img src="images/tit-01.png" style="width:100%" alt="Educación Virtual" />
						<br />
						<p class="btns-v" style="padding-top:10px;text-align:justify;width:75%;margin:0 auto;">
						  	<a href="educacion-virtual.php#educacion-virtual" class="btn btn-danger btn-outline btn-block"  style="">Educación Virtual en la Utec → </a><br>
						  	<a href="educacion-virtual.php#utec-virtual" class="btn btn-danger btn-outline btn-block">UTEC Virtual → </a><br>
						  	<a href="educacion-virtual.php#educacion-exterior" class="btn btn-danger btn-outline btn-block">Educación Virtual en el exterior → </a>
						</p>
						<br />
						<br />
					</div>
				</div>
				<div class="col-ssx-12 col-xs-6 col-sm-8">
					<div class="container-fluid">
						<div class="col-ssx-12 col-xs-6 col-sm-4">
							<a class="black_button" href="http://www.utec.edu.sv/utecvirtualsalvadorenosexterior/" target="_blank">
								<i class="glyphicon glyphicon-info-sign icon-4x"></i><br/> Solicitar Información</a>
							<div class="info_button">Ingresa y conoce un poco mas acerca de las carreras virtuales que ofrece la UTEC.</div>
					    </div>
						<div class="col-ssx-12 col-xs-6 col-sm-4">
							<a class="black_button" href="http://www.utec.edu.sv/utecvirtualsalvadorenosexterior/requisitos/#whatsapplink" target="_blank">
							<i class="glyphicon glyphicon-check icon-4x"></i><br/> Formas de Pago</a>
							<div class="info_button">Descubre las diferentes formas que puedes realizar los pagos de las cuotas de estudio.</div>
						</div>
						<div class="col-ssx-12 col-xs-6 col-sm-4">
							<a class="black_button" href="https://www.utecvirtual.edu.sv/cursos-libres/" target="_blank">
							<i class="glyphicon glyphicon-list-alt icon-4x"></i><br/> Cursos Libres</a>
							<div class="info_button">Aprende mucho mas y conoce nuevas areas a traves de estos cursos mooc.</div>
						</div>
					</div>
				</div>
			</div>
		</div>	
	</section>
	<footer style="background:#343434 url(images/footer-bg.png) bottom repeat-x; padding-top:10px;">
		<div class="container-fluid">
			<div class="row">
				<!-- <div class="col-ssx-12 col-xs-6 col-sm-4" style="text-align:center;color:#fff;"> -->
				 <div class="col-xs-12" style="text-align:center;color:#fff;">
					<h1 style="font-size:1.8em;">UTEC VIRTUAL</h1>
					<p>Universidad Tecnológica de El Salvador<br />
						Calle Arce y 17 Avenida Norte, Edif. José Martí. 2da. Planta, San Salvador, El Salvador, C.A.<br />
						Tels. 2275 - 8723, 2275 - 8888 Ext. 8797
					</p>
				</div>
				<!--
				<div class="col-ssx-12 col-xs-6 col-sm-4 foot-form-solicitud">
					<h2 style="color:#fff;font-size:1.3em;">SOLICITAR INFORMACIÓN</h2>
					<div class="container-fluid">
						<div class="content-form">
							<form id="form1" method="post" action="http://www.utec.edu.sv/distancia/home/post_form/">
								<div class="line">
									<div class="col-xs-6 no-padding">
										<input class="form-control input-sm" type="text" placeholder="Nombres" id="names" name="names">
									</div>
									<div class="col-xs-6 no-padding">
										<input class="form-control input-sm" type="text" placeholder="Apellidos" id="lastnames" name="lastnames">
									</div>
								</div>
								<div class="line">
									<input class="form-control input-sm" type="text" placeholder="Correo electrónico" id="email" name="email">
								</div>
								<div class="line">
									<select class="form-control input-sm" id="carrera" name="carrera">
										<option value="0">Carrera de interés</option>
														<option value="1">Licenciatura en Administración de Empresas</option>
														<option value="2">Licenciatura en Mercadeo</option>
														<option value="3">Ingeniería Industrial</option>
														<option value="4">Ingeniería en Sistemas y Computación</option>
														<option value="5">Licenciatura en Administración de Empresas con Énfasis en Computación</option>
														<option value="6">Licenciatura en Contaduría Pública</option>
														<option value="7">Licenciatura en Informática</option>
									</select>
								</div>
								<div class="line">
									<select onchange="validate_us(this.value);" class="form-control input-sm" id="country" name="pais">
										<option value="0">País</option>
													<option value="75">Estados Unidos</option>
													<option value="42">Canadá</option>
													<option value="1">Afganistán</option>
													<option value="3">Albania</option>
													<option value="4">Alemania</option>
													<option value="5">Andorra</option>
													<option value="6">Angola</option>
													<option value="7">Anguilla</option>
													<option value="8">Antártida</option>
													<option value="9">Antigua y Barbuda</option>
													<option value="10">Antillas Holandesas</option>
													<option value="11">Arabia Saudí</option>
													<option value="12">Argelia</option>
													<option value="13">Argentina</option>
													<option value="14">Armenia</option>
													<option value="15">Aruba</option>
													<option value="131">ARY Macedonia</option>
													<option value="16">Australia</option>
													<option value="17">Austria</option>
													<option value="18">Azerbaiyán</option>
													<option value="19">Bahamas</option>
													<option value="20">Bahréin</option>
													<option value="21">Bangladesh</option>
													<option value="22">Barbados</option>
													<option value="24">Bélgica</option>
													<option value="25">Belice</option>
													<option value="26">Benin</option>
													<option value="27">Bermudas</option>
													<option value="28">Bhután</option>
													<option value="23">Bielorrusia</option>
													<option value="29">Bolivia</option>
													<option value="30">Bosnia y Herzegovina</option>
													<option value="31">Botsuana</option>
													<option value="33">Brasil</option>
													<option value="34">Brunéi</option>
													<option value="35">Bulgaria</option>
													<option value="36">Burkina Faso</option>
													<option value="37">Burundi</option>
													<option value="38">Cabo Verde</option>
													<option value="40">Camboya</option>
													<option value="41">Camerún</option>
													<option value="44">Chad</option>
													<option value="46">Chile</option>
													<option value="47">China</option>
													<option value="48">Chipre</option>
													<option value="50">Ciudad del Vaticano</option>
													<option value="52">Colombia</option>
													<option value="53">Comoras</option>
													<option value="55">Congo</option>
													<option value="57">Corea del Norte</option>
													<option value="58">Corea del Sur</option>
													<option value="59">Costa de Marfil</option>
													<option value="60">Costa Rica</option>
													<option value="61">Croacia</option>
													<option value="62">Cuba</option>
													<option value="63">Dinamarca</option>
													<option value="64">Dominica</option>
													<option value="66">Ecuador</option>
													<option value="67">Egipto</option>
													<option value="68">El Salvador</option>
													<option value="69">Emiratos Árabes Unidos</option>
													<option value="70">Eritrea</option>
													<option value="71">Eslovaquia</option>
													<option value="72">Eslovenia</option>
													<option value="73">España</option>
													<option value="76">Estonia</option>
													<option value="77">Etiopía</option>
													<option value="79">Filipinas</option>
													<option value="80">Finlandia</option>
													<option value="81">Fiyi</option>
													<option value="82">Francia</option>
													<option value="83">Gabón</option>
													<option value="84">Gambia</option>
													<option value="85">Georgia</option>
													<option value="87">Ghana</option>
													<option value="88">Gibraltar</option>
													<option value="89">Granada</option>
													<option value="90">Grecia</option>
													<option value="91">Groenlandia</option>
													<option value="92">Guadalupe</option>
													<option value="93">Guam</option>
													<option value="94">Guatemala</option>
													<option value="95">Guayana Francesa</option>
													<option value="96">Guinea</option>
													<option value="97">Guinea Ecuatorial</option>
													<option value="98">Guinea-Bissau</option>
													<option value="99">Guyana</option>
													<option value="100">Haití</option>
													<option value="102">Honduras</option>
													<option value="103">Hong Kong</option>
													<option value="104">Hungría</option>
													<option value="105">India</option>
													<option value="106">Indonesia</option>
													<option value="107">Irán</option>
													<option value="108">Iraq</option>
													<option value="109">Irlanda</option>
													<option value="32">Isla Bouvet</option>
													<option value="49">Isla de Navidad</option>
													<option value="161">Isla Norfolk</option>
													<option value="110">Islandia</option>
													<option value="39">Islas Caimán</option>
													<option value="51">Islas Cocos</option>
													<option value="56">Islas Cook</option>
													<option value="78">Islas Feroe</option>
													<option value="86">Islas Georgias del Sur y Sandwich del Sur</option>
													<option value="2">Islas Gland</option>
													<option value="101">Islas Heard y McDonald</option>
													<option value="138">Islas Malvinas</option>
													<option value="139">Islas Marianas del Norte</option>
													<option value="141">Islas Marshall</option>
													<option value="174">Islas Pitcairn</option>
													<option value="186">Islas Salomón</option>
													<option value="223">Islas Turcas y Caicos</option>
													<option value="74">Islas ultramarinas de Estados Unidos</option>
													<option value="234">Islas Vírgenes Británicas</option>
													<option value="235">Islas Vírgenes de los Estados Unidos</option>
													<option value="111">Israel</option>
													<option value="112">Italia</option>
													<option value="113">Jamaica</option>
													<option value="114">Japón</option>
													<option value="115">Jordania</option>
													<option value="116">Kazajstán</option>
													<option value="117">Kenia</option>
													<option value="118">Kirguistán</option>
													<option value="119">Kiribati</option>
													<option value="120">Kuwait</option>
													<option value="121">Laos</option>
													<option value="122">Lesotho</option>
													<option value="123">Letonia</option>
													<option value="124">Líbano</option>
													<option value="125">Liberia</option>
													<option value="126">Libia</option>
													<option value="127">Liechtenstein</option>
													<option value="128">Lituania</option>
													<option value="129">Luxemburgo</option>
													<option value="130">Macao</option>
													<option value="132">Madagascar</option>
													<option value="133">Malasia</option>
													<option value="134">Malawi</option>
													<option value="135">Maldivas</option>
													<option value="136">Malí</option>
													<option value="137">Malta</option>
													<option value="140">Marruecos</option>
													<option value="142">Martinica</option>
													<option value="143">Mauricio</option>
													<option value="144">Mauritania</option>
													<option value="145">Mayotte</option>
													<option value="146">México</option>
													<option value="147">Micronesia</option>
													<option value="148">Moldavia</option>
													<option value="149">Mónaco</option>
													<option value="150">Mongolia</option>
													<option value="151">Montserrat</option>
													<option value="152">Mozambique</option>
													<option value="153">Myanmar</option>
													<option value="154">Namibia</option>
													<option value="155">Nauru</option>
													<option value="156">Nepal</option>
													<option value="157">Nicaragua</option>
													<option value="158">Níger</option>
													<option value="159">Nigeria</option>
													<option value="160">Niue</option>
													<option value="162">Noruega</option>
													<option value="163">Nueva Caledonia</option>
													<option value="164">Nueva Zelanda</option>
													<option value="165">Omán</option>
													<option value="166">Países Bajos</option>
													<option value="167">Pakistán</option>
													<option value="168">Palau</option>
													<option value="169">Palestina</option>
													<option value="170">Panamá</option>
													<option value="171">Papúa Nueva Guinea</option>
													<option value="172">Paraguay</option>
													<option value="173">Perú</option>
													<option value="175">Polinesia Francesa</option>
													<option value="176">Polonia</option>
													<option value="177">Portugal</option>
													<option value="178">Puerto Rico</option>
													<option value="179">Qatar</option>
													<option value="180">Reino Unido</option>
													<option value="43">República Centroafricana</option>
													<option value="45">República Checa</option>
													<option value="54">República Democrática del Congo</option>
													<option value="65">República Dominicana</option>
													<option value="181">Reunión</option>
													<option value="182">Ruanda</option>
													<option value="183">Rumania</option>
													<option value="184">Rusia</option>
													<option value="185">Sahara Occidental</option>
													<option value="187">Samoa</option>
													<option value="188">Samoa Americana</option>
													<option value="189">San Cristóbal y Nevis</option>
													<option value="190">San Marino</option>
													<option value="191">San Pedro y Miquelón</option>
													<option value="192">San Vicente y las Granadinas</option>
													<option value="193">Santa Helena</option>
													<option value="194">Santa Lucía</option>
													<option value="195">Santo Tomé y Príncipe</option>
													<option value="196">Senegal</option>
													<option value="197">Serbia y Montenegro</option>
													<option value="198">Seychelles</option>
													<option value="199">Sierra Leona</option>
													<option value="200">Singapur</option>
													<option value="201">Siria</option>
													<option value="202">Somalia</option>
													<option value="203">Sri Lanka</option>
													<option value="204">Suazilandia</option>
													<option value="205">Sudáfrica</option>
													<option value="206">Sudán</option>
													<option value="207">Suecia</option>
													<option value="208">Suiza</option>
													<option value="209">Surinam</option>
													<option value="210">Svalbard y Jan Mayen</option>
													<option value="211">Tailandia</option>
													<option value="212">Taiwán</option>
													<option value="213">Tanzania</option>
													<option value="214">Tayikistán</option>
													<option value="215">Territorio Británico del Océano Índico</option>
													<option value="216">Territorios Australes Franceses</option>
													<option value="217">Timor Oriental</option>
													<option value="218">Togo</option>
													<option value="219">Tokelau</option>
													<option value="220">Tonga</option>
													<option value="221">Trinidad y Tobago</option>
													<option value="222">Túnez</option>
													<option value="224">Turkmenistán</option>
													<option value="225">Turquía</option>
													<option value="226">Tuvalu</option>
													<option value="227">Ucrania</option>
													<option value="228">Uganda</option>
													<option value="229">Uruguay</option>
													<option value="230">Uzbekistán</option>
													<option value="231">Vanuatu</option>
													<option value="232">Venezuela</option>
													<option value="233">Vietnam</option>
													<option value="236">Wallis y Futuna</option>
													<option value="237">Yemen</option>
													<option value="238">Yibuti</option>
													<option value="239">Zambia</option>
													<option value="240">Zimbabue</option>
												</select>
								</div>
								<div class="line">
									<select style="display: none;" class="form-control input-sm"  id="state" name="estado">
										<option value="0">Estado</option>
														<option value="1">Alabama (AL)</option>
														<option value="2">Alaska (AK)</option>
														<option value="3">Arizona (AZ)</option>
														<option value="4">Arkansas (AR)</option>
														<option value="5">California (CA)</option>
														<option value="6">Colorado (CO)</option>
														<option value="7">Connecticut (CT)</option>
														<option value="8">Delaware (DE)</option>
														<option value="9">District of Columbia (DC)</option>
														<option value="10">Florida (FL)</option>
														<option value="11">Georgia (GA)</option>
														<option value="12">Hawaii (HI)</option>
														<option value="13">Idaho (ID)</option>
														<option value="14">Illinois (IL)</option>
														<option value="15">Indiana (IN)</option>
														<option value="16">Iowa (IA)</option>
														<option value="17">Kansas (KS)</option>
														<option value="18">Kentucky (KY)</option>
														<option value="19">Louisiana (LA)</option>
														<option value="20">Maine (ME)</option>
														<option value="21">Maryland (MD)</option>
														<option value="22">Massachusetts (MA)</option>
														<option value="23">Michigan (MI)</option>
														<option value="24">Minnesota (MN)</option>
														<option value="25">Mississippi (MS)</option>
														<option value="26">Missouri (MO)</option>
														<option value="27">Montana (MT)</option>
														<option value="28">Nebraska (NE)</option>
														<option value="29">Nevada (NV)</option>
														<option value="30">New Hampshire (NH)</option>
														<option value="31">New Jersey (NJ)</option>
														<option value="32">New Mexico (NM)</option>
														<option value="33">New York (NY)</option>
														<option value="34">North Carolina (NC)</option>
														<option value="35">North Dakota (ND)</option>
														<option value="36">Ohio (OH)</option>
														<option value="37">Oklahoma (OK)</option>
														<option value="38">Oregon (OR)</option>
														<option value="39">Pennsylvania (PA)</option>
														<option value="40">Rhode Island (RI)</option>
														<option value="41">South Carolina (SC)</option>
														<option value="42">South Dakota (SD)</option>
														<option value="43">Tennessee (TN)</option>
														<option value="44">Texas (TX)</option>
														<option value="45">Utah (UT)</option>
														<option value="46">Vermont (VT)</option>
														<option value="47">Virginia (VA)</option>
														<option value="48">Washington (WA)</option>
														<option value="49">West Virginia (WV)</option>
														<option value="50">Wisconsin (WI)</option>
														<option value="51">Wyoming (WY)</option>
														<option value="52">Ninguno (0)</option>
													</select>
								</div>
								<div class="line">
									<input class="form-control input-sm"  type="text" placeholder="Teléfono" id="tel" name="tel" onkeypress="return validartel(event);">
								</div>
								<div class="line">
								</div>
								<div class="line">
									<input class="form-control input-sm"  type="text" placeholder="Fecha de nacimiento" id="fecha_nac" name="fecha_nac" onkeypress="return false;" onkeyup="return false;" onkeydown="return false" class="hasDatepicker">
								</div>
								<div class="line">
									<select id="medio" name="medio" onchange="show_options(this.value);" class="form-control input-sm">
										<option value="0">¿Por qué medio se enteró?</option>
										<option value="1">Televisión</option>
										<option value="2">Prensa</option>
										<option value="3">Redes sociales</option>
										<option value="4">Web </option>
										<option value="5">Radio</option>
										<option value="7">Visita a Colegios</option>
										<option value="8">Tour Utec</option>
										<option value="6">Otros </option>
									</select>
								</div>
								<div class="line">
									<div id="medio_op1" style="display: none;" class="medios">
										<input type="text" id="canal_medio" name="canal_medio" placeholder="Indique el nombre del canal" class="form-control input-sm" >
									</div>
								</div>
								<div class="line">
									<div id="medio_op2" style="display: none;" class="medios">
										<input type="text" id="periodico_medio" name="periodico_medio" placeholder="Indique el nombre del periódico" class="form-control input-sm" >
									</div>
								</div>
								<div class="line">
									<div id="medio_op3" style="display: none;" class="medios">
										<select id="redsocial" name="redsocial" class="form-control input-sm" >
											<option value="0">Elija la red social</option>
											<option value="Twitter">Twitter</option>
											<option value="Facebook">Facebook</option>
											<option value="Instagram">Instagram</option>
										</select>
								</div>
								</div>
								<div class="line">
									<div id="medio_op4" style="display: none;" class="medios">
										<input type="text" id="web_medio" name="web_medio" placeholder="Indique el nombre o URL del sitio web" class="form-control input-sm" >
									</div>
								</div>
								<div class="line">
									<div id="medio_op5" style="display: none;" class="medios">
										<input type="text" id="radio_medio" name="radio_medio" placeholder="Indique el nombre de la radio" class="form-control input-sm" >
									</div>
								</div>
								<div class="line">
									<div id="medio_op6" style="display: none;" class="medios">
										<input type="text" id="otros_medio" name="otros_medio" placeholder="Indique otro medio" class="form-control input-sm" >
									</div>
								</div>
							</form>
							<img onclick="validate_form();" src="utec/assets/img/bt_enviar.jpg" alt="Enviar">
						</div>
					</div>
					<div id="validatemodal" class="modal hide fade" tabindex="-1" role="dialog" aria-labelledby="myModalLabel" aria-hidden="true">
						<div class="modal-body" id="validatemodal_message"></div>
					</div>

					<div id="yes_modal" class="modal hide fade" tabindex="-1" role="dialog" aria-labelledby="myModalLabel" aria-hidden="true">
					  <div class="modal-body" id="modal_message"> 
						<p>&iexcl;Gracias por completar el formulario, en breve nos comunicaremos con usted!</p>
					  </div>
					</div>
				</div>
				<div class="col-xs-12 col-sm-4" style="text-align:center;">
					
					<img src="images/footer-western.png" style="width:100%" alt="Pagos Via Western Union" />
				</div>
				-->
			</div>
			<div class="row">
				<div style="height:64px;padding:25px">UTEC VIRTUAL &copy;</div>
			</div>
		</div>
	</footer>
	<!-- Area de Mensajes -->
	<div class="modal fade" id="myModal">
	  <div class="modal-dialog" role="document">
		<div class="modal-content">
		  <div class="modal-header">
			<button type="button" class="close" data-dismiss="modal" aria-label="Close">
			  <span aria-hidden="true">&times;</span>
			</button>
			<h4 class="modal-title">Mensaje Importante</h4>
		  </div>
		  <div class="modal-body">
			<p><h4>Estimados alumnos virtuales:</h4><br/>
				Con la finalidad de solventar las dificultades que hemos tenido durante la noche en los servicios virtuales, les notificamos 
				que estarán deshabilitados desde el 23 de  agosto a las 4:00 p.m. hasta el 24 de agosto a las 4:00 p.m.<br/>
				Las evaluaciones y actividades  virtuales de ese periodo serán reprogramadas. 
				Gracias por su comprensión</p>
		  </div>
		  <div class="modal-footer">
			<button type="button" class="btn btn-secondary" data-dismiss="modal">Close</button>
		  </div>
		</div><!-- /.modal-content -->
	  </div><!-- /.modal-dialog -->
	</div><!-- /.modal -->
	<script src="//ajax.googleapis.com/ajax/libs/jquery/1.10.1/jquery.min.js"></script>
    <script>
		window.jQuery || document.write('<script src="js/vendor/jquery-1.10.1.min.js"><\/script>');
		// Obtiene los valores de la fecha, hora, minutos y segundos del servidor
		var jPane = 'time-server';
		var jDate = 'Tuesday, 29 de December del 2015';
		var jHora = '11';
		var jMin = '03';
		var jSec = '50';
		var jTi = 'AM';
	</script>
	<!-- Latest compiled and minified JavaScript -->
	<script src="https://maxcdn.bootstrapcdn.com/bootstrap/3.3.6/js/bootstrap.min.js" integrity="sha384-0mSbJDEHialfmuBBQP6A4Qrprq5OVfW37PRR3j5ELqxss1yVqOtnepnHVP9aJ7xS" crossorigin="anonymous"></script>
	<script src="js/vendor/jssor.slider.mini.js"></script>
	<script src="js/vendor/readmore.min.js"></script>
	<script src="js/vendor/jquery.avgrund.min.js"></script>
	<script src="js/plugins.js?dt=29122017"></script>
    <script src="js/main.js?v1.0.1"></script>
	<script>
		jQuery(document).ready(function ($) {
						//$('#myModal').modal({
			//  show: true
			//});
		
			 var jssor_1_options = {
              $AutoPlay: true,
              $SlideDuration: 4800,
              $Idle: 4000,
              $ArrowKeyNavigation: 0,
              $SlideEasing: $JssorEasing$.$EaseOutQuint,
              $BulletNavigatorOptions: {
                $Class: $JssorBulletNavigator$
              }
            };
            
            var jssor_1_slider = new $JssorSlider$("jssor_1", jssor_1_options);
            
            //responsive code begin
            //you can remove responsive code if you don't want the slider scales while window resizing
            function ScaleSlider() {
                var refSize = jssor_1_slider.$Elmt.parentNode.clientWidth;
                if (refSize) {
                    refSize = Math.min(refSize, 1920);
                    jssor_1_slider.$ScaleWidth(refSize);
                }
                else {
                    window.setTimeout(ScaleSlider, 30);
                }
            }
            ScaleSlider();
            $(window).bind("load", ScaleSlider);
            $(window).bind("resize", ScaleSlider);
            $(window).bind("orientationchange", ScaleSlider);
            //responsive code end


            //Agregamos nuevos elementos a validar
            $("#frmLogin").on('submit',function(e) {
            	var usr = $("#").val(); 
            	var psw = $("#").val(); 
            });

            $(".readmore").readmore({
					speed: 75,
					lessLink: '<a style="text-decoration:none;" href="#">LEER MAS <i class="fa fa-caret-up"></i></a>',
					moreLink: '<a style="text-decoration:none;" href="#">LEER MAS <i class="fa fa-caret-down"></i></a>',
					collapsedHeight: 300,
					embedCSS: false
			});
		});
	</script>
	<script>
	
function validartel(e) 
{
   tecla = e.which || e.keyCode;
   patron = /[0-9\\-]/; // Solo acepta nï¿½meros y guiones
   te = String.fromCharCode(tecla);
   return (patron.test(te) || tecla == 9 || tecla == 8);
}

function validate_us(id)
{
    if(id == 75)
    {
        $("#state").slideDown();
    }
    else
    {
        $("#state").slideUp();
    }
}

function validate_form()
{
    name = $("#names").val();
    apellido = $("#lastnames").val();
    email = $("#email").val();
    carrera = $("#carrera").val();
    pais = $("#country").val();
    estado = $("#state").val();
    tel = $("#tel").val();
    fecha = $("#fecha_nac").val();
    medio = $("#medio").val();
    
    emailPattern = /^[a-zA-Z0-9._-]+@[a-zA-Z0-9.-]+\.[a-zA-Z]{2,4}$/;
    error = "Por favor, corrija los siguientes puntos: <br><br>";
    error_count = 0;
    
    if(name == null || name.length < 2)
    {
        error += " - Escriba su nombre correctamente.<br>";
        error_count++;
    }
    if(apellido == null || apellido.length < 2)
    {
        error += " - Escriba su apellido correctamente.<br>";
        error_count++;
    }
    if(emailPattern.test(email) == false)
    {
        error += " - Digite una direcci&oacute;n de email v&aacute;lida.<br>";
        error_count++;
    }
    if(carrera == 0)
    {
        error += " - Elija la carrera de su inter&eacute;s.<br>";
        error_count++;
    }
    if(pais == 0)
    {
        error += " - Elija su pa&iacute;s de residencia.<br>";
        error_count++;
    }
    if(pais == 75 && estado == 0)
    {
        error += " - Elija su Estado de residencia.<br>";
        error_count++;
    }
    if(tel.length < 7)
    {
        error += " - Indique un n&uacute;mero de tel&eacute;fono v&aacute;lido.<br>";
        error_count++;
    }   
    if(fecha == "")
    {
        error += " - Indique un fecha de nacimiento.<br>";
        error_count++;
    }   
    if(medio == 0)
    {
        error += " - Indique el medio por el cual se enter&oacute;<br>";
        error_count++;
    }
    if(error_count == 0){
        $("#form1").submit();
    }else{
        $("#validatemodal_message").empty();
        $("#validatemodal_message").html(error);
        $("#validatemodal").modal('show');
    }
}

function show_options(opcion)
{
    $("div.medios").slideUp();
    $("div#medio_op" + opcion).slideDown();
}
</script>
<a href="http://www.beyondsecurity.com/vulnerability-scanner-verification/www.utecvirtual.edu.sv"><img src="https://seal.beyondsecurity.com/verification-images/www.utecvirtual.edu.sv/vulnerability-scanner-2.gif" width="0" alt="Website Security Test" border="0" /></a>
</body>
</html>