



<!DOCTYPE html><html lang="es-es"><head><base href="http://www.ujmd.edu.sv/" /><meta http-equiv="content-type" content="text/html; charset=utf-8" /><meta name="keywords" content="universidad, universidades de el salvador, carreras universitarias, ujmd, la matias " /><meta name="robots" content="index, follow" /><meta name="description" content="La Universidad Dr. José Matías Delgado es una corporación de derecho privado, de utilidad pública, sin fines de lucro. " /><title>Universidad Dr. José Matías Delgado | El Salvador - INICIO</title><link href="/?format=feed&amp;type=rss" rel="alternate" type="application/rss+xml" title="RSS 2.0" /><link href="/?format=feed&amp;type=atom" rel="alternate" type="application/atom+xml" title="Atom 1.0" /><link href="/media/com_favicon/icons/1/favicon.ico" rel="shortcut icon" type="image/vnd.microsoft.icon" /><link rel="stylesheet" href="/plugins/system/yt/includes/site/css/style.css" type="text/css" /><link rel="stylesheet" href="http://www.ujmd.edu.sv/media/jbtype/css/font-awesome.css" type="text/css" /><link rel="stylesheet" href="/plugins/system/jcemediabox/css/jcemediabox.css?3ab6d4490e67378d035cce4c84ffa080" type="text/css" /><link rel="stylesheet" href="/plugins/system/jcemediabox/themes/standard/css/style.css?7361405241320e69bc1bfb093eb0a2f7" type="text/css" /><link rel="stylesheet" type="text/css" href="/media/plg_jchoptimize/assets/gz/1/0/aa4a7a1186af0a05211ad43070e9ddd7.css"/><link rel="stylesheet" href="http://fonts.googleapis.com/css?family=Oswald" type="text/css" /><link rel="stylesheet" href="/plugins/system/jabuilder/assets/css/jabuilder.css" type="text/css" /><link rel="stylesheet" href="https://fonts.googleapis.com/icon?family=Material+Icons" type="text/css" /><link rel="stylesheet" href="http://www.ujmd.edu.sv/modules/mod_facebook_slide_likebox/tmpl/css/style1.css" type="text/css" /><link rel="stylesheet" href="/modules/mod_jmnewspro/assets/css/mod_jmnewspro_layout9.css" type="text/css" /><link rel="stylesheet" href="/modules/mod_jmnewspro/assets/css/style_common.css" type="text/css" /><link rel="stylesheet" href="/modules/mod_nice_social_bookmark/css/nsb-opac-inv.css" type="text/css" /><link rel="stylesheet" href="/plugins/content/xtypo/themes/default/style.css" type="text/css" /><link rel="stylesheet" href="/modules/mod_lofarticlesslideshow/assets/jstyle.css" type="text/css" /><style type="text/css">#yt_component .items-leading .item-image{width:540px;max-width:100%;min-height:60px}#yt_component .items-row .item-image{width:210px;max-width:100%;min-height:60px}#yt_menuposition #meganavigator ul.subnavi{position:static;left:auto;right:auto;box-shadow:none}#meganavigator ul.subnavi>li{margin-left:0}#meganavigator ul.subnavi>li.first{margin-top:0}body.sj_news{font-size:12px}body.sj_news{font-family:arial,sans-serif}.google-font,.modtitle,li.level1>.item-link,div.mega-group-title,.related-items-title,.page-header h1,h1.heading-category,div.pagination ul.pagination{font-family:Oswald,serif !important}body.sj_news{background-color:#fff;color:#000}body a{color:#00f}#yt_header{background-color:#100159}#yt_spotlight3{background-color:#242963}#yt_spotlight4{background-color:#00487c}#yt_footer{background-color:#0f0f0f}#yt_spotlight5{background-color:#00487c}#jmnewspro-151 .bx-pager{display:none}#jmnewspro-151 .bx-controls{left:0;position:absolute;bottom:-15px}.nsb_container a.icons{padding:px;float:left;display:inline-block}#plusone{padding:px !important}#goog-gt-tt{display:none !important}.goog-te-banner-frame{display:none !important}.goog-te-menu-value:hover{text-decoration:none !important}body{top:0 !important}#google_translate_element2{display:none!important}a.flag{font-size:24px;padding:1px 0;background-repeat:no-repeat;background-image:url('/modules/mod_gtranslate/tmpl/lang/24a.png')}a.flag:hover{background-image:url('/modules/mod_gtranslate/tmpl/lang/24.png')}a.flag img{border:0}a.alt_flag{font-size:24px;padding:1px 0;background-repeat:no-repeat;background-image:url('/modules/mod_gtranslate/tmpl/lang/alt_flagsa.png')}a.alt_flag:hover{background-image:url('/modules/mod_gtranslate/tmpl/lang/alt_flags.png')}a.alt_flag img{border:0}</style> <script src="/plugins/system/yt/includes/admin/js/jquery.min.js" type="text/javascript"></script> <script src="/plugins/system/yt/includes/admin/js/jquery-noconflict.js" type="text/javascript"></script> <script src="/media/jui/js/jquery.min.js" type="text/javascript"></script> <script type="application/javascript" src="/media/plg_jchoptimize/assets/gz/1/0/5883126907234e5810d2b828660b554b.js"></script> <script src="/media/jui/js/jquery-migrate.min.js" type="text/javascript"></script> <script type="application/javascript" src="/media/plg_jchoptimize/assets/gz/1/1/5883126907234e5810d2b828660b554b.js"></script> <script src="/plugins/system/jcemediabox/js/jcemediabox.js?2ee2100a9127451a41de5a4c2c62e127" type="text/javascript"></script> <script type="application/javascript" src="/media/plg_jchoptimize/assets/gz/1/2/5883126907234e5810d2b828660b554b.js"></script> <script src="/plugins/system/jabuilder/assets/js/jabuilder.js" type="text/javascript"></script> <script src="/modules/mod_jmnewspro/assets/js/jquery.bxslider.js" type="text/javascript"></script> <script src="/modules/mod_jmnewspro/assets/js/jquery.easing.1.3.js" type="text/javascript"></script> <script src="/modules/mod_jmnewspro/assets/js/jquery.jm-bxslider.js" type="text/javascript"></script> <script src="/plugins/content/xtypo/assets/script.js" type="text/javascript"></script> <script type="application/javascript" src="/media/plg_jchoptimize/assets/gz/1/3/5883126907234e5810d2b828660b554b.js"></script> <script src="/modules/mod_lofarticlesslideshow/assets/jscript.js" type="text/javascript"></script> <script type="text/javascript">jQuery(window).on('load',function(){new JCaption('img.caption');});JCEMediaBox.init({popup:{width:"",height:"",legacy:0,lightbox:0,shadowbox:0,resize:1,icons:1,overlay:1,overlayopacity:0.8,overlaycolor:"#000000",fadespeed:500,scalespeed:500,hideobjects:0,scrolling:"fixed",close:2,labels:{'close':'Cerrar','next':'Siguiente','previous':'Anterior','cancel':'Cancelar','numbers':'{$current} de {$total}'},cookie_expiry:"",google_viewer:0},tooltip:{className:"tooltip",opacity:0.8,speed:150,position:"br",offsets:{x:16,y:16}},base:"/",imgpath:"plugins/system/jcemediabox/img",theme:"standard",themecustom:"",themepath:"plugins/system/jcemediabox/themes",mediafallback:0,mediaselector:"audio,video"});function responsiveTables(){for(var e=document.querySelectorAll("table"),t=0;t<e.length;t++)if(e[t].scrollWidth>e[t].parentNode.clientWidth&&("div"!=e[t].parentNode.tagName.toLowerCase()||"res-div"!=e[t].parentNode.getAttribute("data-responsive"))){var r=document.createElement("div"),o=e[t].parentNode;r.appendChild(document.createTextNode("Desplácese hacia la derecha para obtener más ->")),r.appendChild(e[t].cloneNode(!0)),r.setAttribute("style","overflow-x:scroll;"),r.setAttribute("data-responsive","res-div"),o.replaceChild(r,e[t])}else if(e[t].scrollWidth<=e[t].parentNode.clientWidth&&"div"==e[t].parentNode.tagName.toLowerCase()&&"res-div"==e[t].parentNode.getAttribute("data-responsive")){var a=e[t].parentNode,d=a.parentNode;d.replaceChild(e[t].cloneNode(!0),a)}}window.addEventListener("resize",function(){responsiveTables()}),document.onreadystatechange=function(){"complete"==document.readyState&&responsiveTables()};(function(d){var js,id='powr-js',ref=d.getElementsByTagName('script')[0];if(d.getElementById(id)){return;}
js=d.createElement('script');js.id=id;js.async=true;js.src='http://www.ujmd.edu.sv/plugins/content/powrshortcodes/powr_joomla.js';js.setAttribute('powr-token','j6qOADUkbU1491514895');js.setAttribute('external-type','joomla');ref.parentNode.insertBefore(js,ref);}(document));(function(d){var js,id='powr-js',ref=d.getElementsByTagName('script')[0];if(d.getElementById(id)){return;}
js=d.createElement('script');js.id=id;js.async=true;js.src='http://www.ujmd.edu.sv/plugins/content/powrshortcodes/powr_joomla.js';js.setAttribute('powr-token','j6qOADUkbU1491514895');js.setAttribute('external-type','joomla');ref.parentNode.insertBefore(js,ref);}(document));</script> <script type="text/javascript">var TMPL_NAME="sj_news";var TMPL_COOKIE=["direction","fontSize","fontName","templateColor","bgcolor","linkcolor","textcolor","header-bgimage","header-bgcolor","spotlight3-bgcolor","spotlight4-bgcolor","spotlight5-bgcolor","footer-bgcolor","footer-bgimage","templateLayout","menustyle","googleWebFont","activeNotice"];function MobileRedirectUrl(){window.location.href=document.getElementById("yt-mobilemenu").value;}</script> <script type="text/javascript">window.addEvent("domready",function(){if(typeof jQuery!="undefined"&&typeof MooTools!="undefined"){Element.implement({hide:function(how,mode){return this;}});}});</script> <script type="text/javascript" src="http://s7.addthis.com/js/300/addthis_widget.js"></script><meta name="HandheldFriendly" content="true"/><meta name="viewport" content="width=device-width, target-densitydpi=160dpi, minimum-scale=1.0, maximum-scale=1.0, user-scalable=no" /><meta http-equiv="content-type" content="text/html; charset=utf-8" /><!--[ if lt IE 9]>
<script src="http://www.ujmd.edu.sv/templates/sj_news/js/respond.min.js" type="text/javascript"></script>
<script src="http://www.ujmd.edu.sv/templates/sj_news/js/modernizr.min.js" type="text/javascript"></script>
<script src="http://html5shiv.googlecode.com/svn/trunk/html5.js"> </ script>
<[endif] --> <!--For param enableGoogleAnalytics--> <script type="text/javascript">var _gaq=_gaq||[];_gaq.push(["_setAccount","UA-42640012-1"]);_gaq.push(["_trackPageview"]);(function(){var ga=document.createElement("script");ga.type="text/javascript";ga.async=true;ga.src=("https:"==document.location.protocol?"https://ssl":"http://www")+".google-analytics.com/ga.js";var s=document.getElementsByTagName("script")[0];s.parentNode.insertBefore(ga,s);})();</script> <!-- Facebook Pixel Code --> <script>!function(f,b,e,v,n,t,s){if(f.fbq)return;n=f.fbq=function(){n.callMethod?n.callMethod.apply(n,arguments):n.queue.push(arguments)};if(!f._fbq)f._fbq=n;n.push=n;n.loaded=!0;n.version='2.0';n.queue=[];t=b.createElement(e);t.async=!0;t.src=v;s=b.getElementsByTagName(e)[0];s.parentNode.insertBefore(t,s)}(window,document,'script','https://connect.facebook.net/en_US/fbevents.js');fbq('init','155114058295102');fbq('track','PageView');</script><noscript><img height="1" width="1" style="display:none"
src="https://www.facebook.com/tr?id=155114058295102&ev=PageView&noscript=1"
/></noscript><!-- DO NOT MODIFY --> <!-- End Facebook Pixel Code --> <script>(function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){(i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)})(window,document,'script','//www.google-analytics.com/analytics.js','ga');ga('create','UA-113032910-1','http://www.ujmd.edu.sv');ga('send','pageview');</script> <!-- Universal Google Analytics Plugin by PB Web Development --> </head><body id="bd" class="homepage com_content view-featured blue sj_news layout_main-right.xml no-slideshow  yt-jv3" onLoad="prettyPrint()"><style type="text/css">body{background-image:url("http://www.ujmd.edu.sv/images/Fotos_para_Contenido/Fondo_Sitio_Web_blanco2.jpg")!important;background-attachment:fixed!important;background-position:center center!important;background-repeat:repeat!important;background-color:transparent!important}</style><section id="yt_wrapper"> <a id="top" name="scroll-to-top"></a> <header id="yt_header" class="block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="yt_logoposition" class="span3" data-normal="span3" data-tablet="span3" data-stablet="span3"> <a href="/index.php" title="Universidad Dr. José Matías Delgado | El Salvador"> <img alt="Universidad Dr. José Matías Delgado | El Salvador" src="http://www.ujmd.edu.sv/images/logoujmdv2.png"/> </a> </div><div id="position-0" class="span5 offset4" data-normal="span5 offset4" data-tablet="span5 offset4" data-stablet="span7 offset2"><div id="yt_searchcustom"> <a class="btn-seach"></a> <form action="/" method="post"><div class="search"> <!--<label for="mod-search-searchword">Buscar...</label>--><input name="searchword" id="mod_search_searchword" maxlength="200" alt="Buscar" class="inputbox" type="text" size="20" value="Buscar..." onblur="if(this.value=='') this.value='Buscar...';" onfocus="if(this.value=='Buscar...') this.value='';" /><input type="submit" value="Buscar" class="button" onclick="this.form.searchword.focus();"/> <input type="hidden" name="task" value="search" /> <input type="hidden" name="option" value="com_search" /> <input type="hidden" name="Itemid" value="101" /> </div></form></div><noscript>Javascript is required to use <a href="http://gtranslate.net/">GTranslate</a> <a href="http://gtranslate.net/">multilingual website</a> and <a href="http://gtranslate.net/">translation delivery network</a></noscript> <script type="text/javascript">eval(function(p,a,c,k,e,r){e=function(c){return(c<a?'':e(parseInt(c/a)))+((c=c%a)>35?String.fromCharCode(c+29):c.toString(36))};if(!''.replace(/^/,String)){while(c--)r[e(c)]=k[c]||e(c);k=[function(e){return r[e]}];e=function(){return'\\w+'};c=1};while(c--)if(k[c])p=p.replace(new RegExp('\\b'+e(c)+'\\b','g'),k[c]);return p}('6 7(a,b){n{4(2.9){3 c=2.9("o");c.p(b,f,f);a.q(c)}g{3 c=2.r();a.s(\'t\'+b,c)}}u(e){}}6 h(a){4(a.8)a=a.8;4(a==\'\')v;3 b=a.w(\'|\')[1];3 c;3 d=2.x(\'y\');z(3 i=0;i<d.5;i++)4(d[i].A==\'B-C-D\')c=d[i];4(2.j(\'k\')==E||2.j(\'k\').l.5==0||c.5==0||c.l.5==0){F(6(){h(a)},G)}g{c.8=b;7(c,\'m\');7(c,\'m\')}}',43,43,'||document|var|if|length|function|GTranslateFireEvent|value|createEvent||||||true|else|doGTranslate||getElementById|google_translate_element2|innerHTML|change|try|HTMLEvents|initEvent|dispatchEvent|createEventObject|fireEvent|on|catch|return|split|getElementsByTagName|select|for|className|goog|te|combo|null|setTimeout|500'.split('|'),0,{}))</script><div id="google_translate_element2"></div> <script type="text/javascript">function googleTranslateElementInit2(){new google.translate.TranslateElement({pageLanguage:'es',autoDisplay:false},'google_translate_element2');}</script> <script type="text/javascript" src="http://translate.google.com/translate_a/element.js?cb=googleTranslateElementInit2"></script> <a href="#" onclick="doGTranslate('es|es');return false;" title="Spanish" class="flag nturl" style="background-position:-600px -200px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="24" width="24" alt="Spanish" /></a> <a href="#" onclick="doGTranslate('es|en');return false;" title="English" class="alt_flag" style="background-position:-0px -100px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="24" width="24" alt="English" /></a> <a href="#" onclick="doGTranslate('es|fr');return false;" title="French" class="flag nturl" style="background-position:-200px -100px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="24" width="24" alt="French" /></a> <a href="#" onclick="doGTranslate('es|it');return false;" title="Italian" class="flag nturl" style="background-position:-600px -100px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="24" width="24" alt="Italian" /></a> </div></div></div></div></header><section id="yt_menuwrap" class="block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="yt_menuposition" class="span12"><ul id="meganavigator" class="navi"><li class="active level1 first"> <a class="active level1 first item-link" href="http://www.ujmd.edu.sv/"><span class="menu-title">INICIO</span></a> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">LA UNIVERSIDAD </span></div><!-- open mega-content div --><div class="level2 mega-content" ><div class="mega-content-inner" style="width:400px"><div class="mega-col first more" style="width:200px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/la-universidad/institución"><span class="menu-title">Institución</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/la-universidad/campus"><span class="menu-title">Ubicación de Unidades Académicas y Administrativas</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/la-universidad/acreditación-y-convenios"><span class="menu-title">Acreditación, Certificación y Convenios </span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/la-universidad/unidades-de-apoyo-académico-administrativas"><span class="menu-title">Unidades Académico-administrativas </span></a> </li> </ul> </div><div class="mega-col last more" style="width:200px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/la-universidad/incorporaciones"><span class="menu-title">Incorporaciones</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/la-universidad/todas-las-noticias"><span class="menu-title">Noticias Archivadas </span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/la-universidad/especial-40-anos"><span class="menu-title">Especial 40 años</span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">ADMISIÓN</span></div><div class="level2 mega-content" ><div class="mega-content-inner" ><div class="mega-col first one" ><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/admisión/nuevo-ingreso-e-ingreso-por-equivalencia"><span class="menu-title">Nuevo Ingreso e Ingreso por Equivalencia </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/admisión/proceso-de-reingreso"><span class="menu-title">Proceso de Reingreso </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/admisión/horarios-cursillo-preuniversitario"><span class="menu-title">Horarios Cursillo Preuniversitario</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/admisión/resultados-del-cursillo-pre-universitario"><span class="menu-title">Resultados del Cursillo Pre-universitario </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/admisión/aranceles"><span class="menu-title">Aranceles </span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/admisión/becas"><span class="menu-title">Becas </span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">OFERTA ACADÉMICA</span></div><div class="level2 mega-content" ><div class="mega-content-inner" ><div class="mega-col first one" ><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/oferta-académica/facultades-y-escuelas"><span class="menu-title">Facultades </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/oferta-académica/carreras-universitarias"><span class="menu-title">Carreras Universitarias </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/oferta-académica/programas-de-posgrado"><span class="menu-title">Posgrados y Educación Continua</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/oferta-académica/centro-de-idiomas"><span class="menu-title">Centro de idiomas</span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="http://matiasvirtual.net" target="_blank"><span class="menu-title">Aulas virtuales</span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">CICLO ACADÉMICO </span></div><div class="level2 mega-content" ><div class="mega-content-inner" style="width:500px"><div class="mega-col first more" style="width:250px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/ciclo-académico/calendario-académico"><span class="menu-title">Calendario Académico </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/ciclo-académico/horarios-de-inscripción"><span class="menu-title">Horarios de Inscripción </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/ciclo-académico/horarios-de-clases"><span class="menu-title">Horarios de Clases</span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/ciclo-académico/horarios-de-parciales"><span class="menu-title">Horarios de Parciales </span></a> </li> </ul> </div><div class="mega-col last more" style="width:250px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/ciclo-académico/horarios-de-seminarios-de-investigación-y-especialización"><span class="menu-title">Horarios de Seminarios de Investigación y Especialización</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/ciclo-académico/cursos-de-formación-complementaria"><span class="menu-title">Cursos de Formación Complementarias</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/ciclo-académico/ofertas-para-servicio-social"><span class="menu-title">Ofertas para Servicio Social</span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/ciclo-académico/facultad-de-economía,-empresa-y-negocios-proceso-de-graduación"><span class="menu-title">Facultad de Economía, Empresa y Negocios: Proceso de Graduación</span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">SERVICIOS </span></div><div class="level2 mega-content" ><div class="mega-content-inner" style="width:500px"><div class="mega-col first more" style="width:250px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/servicios-universitarios/servicios-de-la-universidad"><span class="menu-title">Servicios de la Universidad </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/servicios-universitarios/servicios-en-línea"><span class="menu-title">Servicios en Línea</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/servicios-universitarios/imagen-institucional"><span class="menu-title">Formularios de Imagen Institucional </span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/servicios-universitarios/bolsa-de-trabajo-ujmd"><span class="menu-title">Bolsa de Trabajo UJMD </span></a> </li> </ul> </div><div class="mega-col last more" style="width:250px;"><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/servicios-universitarios/mapa-del-sitio"><span class="menu-title">Mapa del sitio</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/servicios-universitarios/directorio-telefonico-ujmd"><span class="menu-title">Directorio Telefónico UJMD</span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/servicios-universitarios/clinica-matias"><span class="menu-title">Clínica de Asistencia Psicológica</span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">INVESTIGACIÓN</span></div><div class="level2 mega-content" ><div class="mega-content-inner" ><div class="mega-col first one" ><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="http://cich.ujmd.edu.sv" target="_blank"><span class="menu-title">Centro de Investigaciones en Ciencias y Humanidades (CICH)</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/investigación/revistas-digitales"><span class="menu-title">Revistas Digitales </span></a> </li> <li class="level2"> <a class="level2 item-link" href="http://iij.ujmd.edu.sv/" target="_blank"><span class="menu-title">Instituto de Investigación Jurídica IIJ</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/investigación/investigaciones-de-posgrados"><span class="menu-title">Investigaciones de Posgrados</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/investigación/editorial-delgado-stand-virtual"><span class="menu-title">Editorial Delgado Stand Virtual</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/investigación/observatorio-virtual"><span class="menu-title">Observatorio Virtual</span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/investigación/comite-de-etica-de-la-investigacion-en-salud-ujmd-ceis-ujmd"><span class="menu-title">Comité de Ética de la Investigación en Salud- UJMD (CEIS-UJMD)</span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 havechild"><div class="level1 havechild item-link separator"><span class="menu-title">Proyección Social</span></div><div class="level2 mega-content" ><div class="mega-content-inner" ><div class="mega-col first one" ><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="/proyeccion-social/proyectos-desarrollados"><span class="menu-title">Proyectos Desarrollados </span></a> </li> </ul> </div> </div> </div> </li> <li class="level1 last havechild"><div class="level1 last havechild item-link separator"><span class="menu-title">Docencia</span></div><div class="level2 mega-content" ><div class="mega-content-inner" ><div class="mega-col first one" ><ul class="subnavi level2"><li class="level2 first"> <a class="level2 first item-link" href="https://www.google.com/url?q=https%3A%2F%2Fdevujmd.wixsite.com%2Fpdecap2018dev&amp;sa=D&amp;sntz=1&amp;usg=AFQjCNF2uwFJC8IMbmqWzcAPjztzt_1Yww"><span class="menu-title">Programas de Capacitación</span></a> </li> <li class="level2"> <a class="level2 item-link" href="/docencia/dirección-de-informática"><span class="menu-title">Dirección de Informática </span></a> </li> <li class="level2"> <a class="level2 item-link" href="/docencia/desarrollo-y-seguimiento-curricular"><span class="menu-title">Desarrollo y Seguimiento Curricular</span></a> </li> <li class="level2"> <a class="level2 item-link" href="https://accounts.google.com/ServiceLogin?service=mail&amp;continue=https://mail.google.com/mail/&amp;hl=es" target="_blank"><span class="menu-title">Correo Institucional </span></a> </li> <li class="level2 last"> <a class="level2 last item-link" href="/docencia/dirección-de-educación-virtual"><span class="menu-title">Dirección de Educación Virtual</span></a> </li> </ul> </div> </div> </div> </li> </ul> <script type="text/javascript">jQuery(function($){$('#meganavigator').megamenu({'wrap':'#yt_menuwrap .container','easing':'easeOutCirc','speed':'500','justify':'left'});});</script> <select id="yt-mobilemenu" name="menu" onchange="MobileRedirectUrl()"> <option selected="selected" value='http://www.ujmd.edu.sv/'>INICIO</option> <option value="#1">LA UNIVERSIDAD </option> <option value='/la-universidad/institución'>-- Institución</option> <option value='/la-universidad/campus'>-- Ubicación de Unidades Académicas y Administrativas</option> <option value='/la-universidad/acreditación-y-convenios'>-- Acreditación, Certificación y Convenios </option> <option value='/la-universidad/unidades-de-apoyo-académico-administrativas'>-- Unidades Académico-administrativas </option> <option value='/la-universidad/incorporaciones'>-- Incorporaciones</option> <option value='/la-universidad/todas-las-noticias'>-- Noticias Archivadas </option> <option value='/la-universidad/especial-40-anos'>-- Especial 40 años</option> <option value="#1">ADMISIÓN</option> <option value='/admisión/nuevo-ingreso-e-ingreso-por-equivalencia'>-- Nuevo Ingreso e Ingreso por Equivalencia </option> <option value='/admisión/proceso-de-reingreso'>-- Proceso de Reingreso </option> <option value='/admisión/horarios-cursillo-preuniversitario'>-- Horarios Cursillo Preuniversitario</option> <option value='/admisión/resultados-del-cursillo-pre-universitario'>-- Resultados del Cursillo Pre-universitario </option> <option value='/admisión/aranceles'>-- Aranceles </option> <option value='/admisión/becas'>-- Becas </option> <option value="#1">OFERTA ACADÉMICA</option> <option value='/oferta-académica/facultades-y-escuelas'>-- Facultades </option> <option value='/oferta-académica/carreras-universitarias'>-- Carreras Universitarias </option> <option value='/oferta-académica/programas-de-posgrado'>-- Posgrados y Educación Continua</option> <option value='/oferta-académica/centro-de-idiomas'>-- Centro de idiomas</option> <option value='http://matiasvirtual.net'>-- Aulas virtuales</option> <option value="#1">CICLO ACADÉMICO </option> <option value='/ciclo-académico/calendario-académico'>-- Calendario Académico </option> <option value='/ciclo-académico/horarios-de-inscripción'>-- Horarios de Inscripción </option> <option value='/ciclo-académico/horarios-de-clases'>-- Horarios de Clases</option> <option value='/ciclo-académico/horarios-de-parciales'>-- Horarios de Parciales </option> <option value='/ciclo-académico/horarios-de-seminarios-de-investigación-y-especialización'>-- Horarios de Seminarios de Investigación y Especialización</option> <option value='/ciclo-académico/cursos-de-formación-complementaria'>-- Cursos de Formación Complementarias</option> <option value='/ciclo-académico/ofertas-para-servicio-social'>-- Ofertas para Servicio Social</option> <option value='/ciclo-académico/facultad-de-economía,-empresa-y-negocios-proceso-de-graduación'>-- Facultad de Economía, Empresa y Negocios: Proceso de Graduación</option> <option value="#1">SERVICIOS </option> <option value='/servicios-universitarios/servicios-de-la-universidad'>-- Servicios de la Universidad </option> <option value='/servicios-universitarios/servicios-en-línea'>-- Servicios en Línea</option> <option value='/servicios-universitarios/imagen-institucional'>-- Formularios de Imagen Institucional </option> <option value='/servicios-universitarios/bolsa-de-trabajo-ujmd'>-- Bolsa de Trabajo UJMD </option> <option value='/servicios-universitarios/mapa-del-sitio'>-- Mapa del sitio</option> <option value='/servicios-universitarios/directorio-telefonico-ujmd'>-- Directorio Telefónico UJMD</option> <option value='/servicios-universitarios/clinica-matias'>-- Clínica de Asistencia Psicológica</option> <option value="#1">INVESTIGACIÓN</option> <option value='http://cich.ujmd.edu.sv'>-- Centro de Investigaciones en Ciencias y Humanidades (CICH)</option> <option value='/investigación/revistas-digitales'>-- Revistas Digitales </option> <option value='http://iij.ujmd.edu.sv/'>-- Instituto de Investigación Jurídica IIJ</option> <option value='/investigación/investigaciones-de-posgrados'>-- Investigaciones de Posgrados</option> <option value='/investigación/editorial-delgado-stand-virtual'>-- Editorial Delgado Stand Virtual</option> <option value='/investigación/observatorio-virtual'>-- Observatorio Virtual</option> <option value='/investigación/comite-de-etica-de-la-investigacion-en-salud-ujmd-ceis-ujmd'>-- Comité de Ética de la Investigación en Salud- UJMD (CEIS-UJMD)</option> <option value="#1">Proyección Social</option> <option value='/proyeccion-social/proyectos-desarrollados'>-- Proyectos Desarrollados </option> <option value="#1">Docencia</option> <option value='https://www.google.com/url?q=https%3A%2F%2Fdevujmd.wixsite.com%2Fpdecap2018dev&amp;sa=D&amp;sntz=1&amp;usg=AFQjCNF2uwFJC8IMbmqWzcAPjztzt_1Yww'>-- Programas de Capacitación</option> <option value='/docencia/dirección-de-informática'>-- Dirección de Informática </option> <option value='/docencia/desarrollo-y-seguimiento-curricular'>-- Desarrollo y Seguimiento Curricular</option> <option value='https://accounts.google.com/ServiceLogin?service=mail&amp;continue=https://mail.google.com/mail/&amp;hl=es'>-- Correo Institucional </option> <option value='/docencia/dirección-de-educación-virtual'>-- Dirección de Educación Virtual</option> </select> </div></div></div></div></section><section id="yt_slideshow" class="block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="slideshow" class="span8" data-normal="" data-tablet="" data-stablet="span12"><div class="module "><div class="modcontent clearfix"><div id="lofass156" class="lof-ass " style="height:auto; width:auto"><div class="lofass-container  lof-css3  "><div class="preload"><div></div></div><div class="lof-main-wapper" style="height:350px;width:620px;"><div class="lof-main-item "> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-gradvirting.png" title="Graduación Virtual Facultad de Ingeniería" width="620" alt="Graduación Virtual Facultad de Ingeniería" > <div class="lof-description"><h4><a target="_parent" title="Graduación Virtual Facultad de Ingeniería" href="/contenidoslideshow/29-noticias/2182-graduacion-virtual-facultad-de-ingenieria-2">Graduación Virtual Facultad de Ingeniería</a></h4><p>Este viernes 16 de marzo de 2018 se llev&oacute; a cabo una Graduaci&oacute;n Virtual por parte de la Facultad de Ingenier&iacute;a, en las...</p></div></div><div class="lof-main-item"> <img src="/images/Redacci&oacute;nMultimedia.png" title="ECC: Evaluación de trabajos periodísticos multimedia" width="620" alt="ECC: Evaluación de trabajos periodísticos multimedia" > <div class="lof-description"><h4><a target="_parent" title="ECC: Evaluación de trabajos periodísticos multimedia" href="/contenidoslideshow/29-noticias/2181-ecc-evaluacion-de-trabajos-periodisticos-multimedia">ECC: Evaluación de trabajos periodísticos multimedia</a></h4><p>El pasado viernes 16 de marzo, los estudiantes de la c&aacute;tedra G&eacute;neros Period&iacute;sticos, (materia optativa), impartida por el...</p></div></div><div class="lof-main-item"> <img src="/images/Afiche_ABC_del_&eacute;xito_empresarial-1.jpg" title="Expertos del TEC impartirán Diplomado "ABC del Éxito Empresarial"" width="620" alt="Expertos del TEC impartirán Diplomado "ABC del Éxito Empresarial"" > <div class="lof-description"><h4><a target="_parent" title="Expertos del TEC impartirán Diplomado "ABC del Éxito Empresarial"" href="/contenidoslideshow/29-noticias/2180-expertos-del-tec-impartiran-diplomado-abc-del-exito-empresarial">Expertos del TEC impartirán Diplomado "ABC del Éxito Empresarial"</a></h4><p> &nbsp; </p></div></div><div class="lof-main-item"> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-yomeSumocintillo.jpg" title="Invitación a la presentación de los resultados del proyecto #YoMeSumo" width="620" alt="Invitación a la presentación de los resultados del proyecto #YoMeSumo" > <div class="lof-description"><h4><a target="_parent" title="Invitación a la presentación de los resultados del proyecto #YoMeSumo" href="/contenidoslideshow/29-noticias/2178-invitacion-a-la-presentacion-de-los-resultados-del-proyecto-yomesumo">Invitación a la presentación de los resultados del proyecto #YoMeSumo</a></h4><p>Comunidad Mat&iacute;as te invitamos a participar en el evento: </p></div></div><div class="lof-main-item"> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-evaluarnoticias.png" title="Completa la "Evaluación Docente"" width="620" alt="Completa la "Evaluación Docente"" > <div class="lof-description"><h4><a target="_parent" title="Completa la "Evaluación Docente"" href="/contenidoslideshow/29-noticias/2156-completa-la-evaluacion-docente">Completa la "Evaluación Docente"</a></h4><p>Estimado estudiante te notificamos que ya puedes completar la "Evaluaci&oacute;n Docente", tu participaci&oacute;n es clave para mejorar la...</p></div></div><div class="lof-main-item"> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-derechoprivados.JPG" title="Privados escritos abril 2018" width="620" alt="Privados escritos abril 2018" > <div class="lof-description"><h4><a target="_parent" title="Privados escritos abril 2018" href="/contenidoslideshow/29-noticias/2104-privados-escritos-abril-2018">Privados escritos abril 2018</a></h4><p></p></div></div><div class="lof-main-item"> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-hugolindoportada.png" title="Participa en Premio Hugo Lindo de Novela" width="620" alt="Participa en Premio Hugo Lindo de Novela" > <div class="lof-description"><h4><a target="_parent" title="Participa en Premio Hugo Lindo de Novela" href="/contenidoslideshow/29-noticias/2041-participa-en-premio-hugo-lindo-de-novela">Participa en Premio Hugo Lindo de Novela</a></h4><p>Editorial Delgado te invita a participar en el Premio Hugo Lindo de Novela 2018 Como parte del 40 aniversario de fundaci&oacute;n, la universidad...</p></div></div><div class="lof-main-item"> <img src="http://www.ujmd.edu.sv/cache/lofthumbs/620x350-capacitaciondocente.png" title="Programa de Capacitación en línea para personal Docente y Administrativo" width="620" alt="Programa de Capacitación en línea para personal Docente y Administrativo" > <div class="lof-description"><h4><a target="_parent" title="Programa de Capacitación en línea para personal Docente y Administrativo" href="/contenidoslideshow/29-noticias/1896-programa-de-capacitacion-en-linea-para-personal-docente-y-administrativo">Programa de Capacitación en línea para personal Docente y Administrativo</a></h4><p>Comunidad Mat&iacute;as: La Facultad de Posgrados y Educaci&oacute;n Continua,&nbsp;Direcci&oacute;n de Recursos Humanos y&nbsp;la...</p></div></div></div><div class="lof-buttons-control"> <a href="/" onclick="return false;" class="lof-previous">Previous</a> <a href="/" class="lof-next" onclick="return false;">Next</a> </div></div></div> <script type="text/javascript">var _lofmain=$('lofass156');var object=new LofArticleSlideshow(_lofmain,{fxObject:{transition:Fx.Transitions.Quad.easeInOut,duration:500},startItem:0,interval:5000,direction:'hrleft',navItemHeight:100,navItemWidth:310,navItemsDisplay:3,navPos:'0',autoStart:1,descOpacity:1});object.registerButtonsControl('click',{next:_lofmain.getElement('.lof-next'),previous:_lofmain.getElement('.lof-previous')});</script> </div> </div> </div><div id="position-1" class="span4" data-normal="" data-tablet="" data-stablet="span12 first"><div class="module "><h3 class="modtitle">Síguenos en:</h3><div class="modcontent clearfix"><div class="nsb_container"><a id="l1" class="icons" target="_blank" href="http://www.facebook.com/UniversidadDrJoseMatiasDelgado"><img title="Facebook" src="/modules/mod_nice_social_bookmark/icons/facebook_aqu_32.png" alt="Facebook" /></a><a id="l3" class="icons" target="_blank" href="http://www.twitter.com/#!/UJMD_sv"><img title="Twitter" src="/modules/mod_nice_social_bookmark/icons/twitter_aqu_32.png" alt="Twitter" /></a><a id="ll1" class="icons" target="_blank" href="http://www.linkedin.com/in/ujmd-mat%C3%ADas-delgado/"><img title="LinkedIn" src="/modules/mod_nice_social_bookmark/icons/linkedin_aqu_32.png" alt="LinkedIn" /></a><a id="l21" class="icons" target="_blank" href="http://pinterest.com/ujmd"><img title="Pinterest" src="/modules/mod_nice_social_bookmark/icons/pinterest_aqu_32.png" alt="Pinterest" /></a><a id="l16" class="icons" target="_blank" href="http://www.youtube.com/user/MatiasUJMD"><img title="" src="/images/Fotos_para_Contenido/youtube-2-icon.png" alt="YouTube" /></a><a id="l17" class="icons" target="_blank" href="https://plus.google.com/u/0/+UjmdEduSvUJMD/posts"><img title="" src="/images/Fotos_para_Contenido/Google_plus.png" alt="Google+" /></a><a id="l18" class="icons" target="_blank" href="https://www.instagram.com/universidad_ujmd/"><img title="" src="/images/Fotos_para_Contenido/Instagram.png" alt="Instagram" /></a></div><div style="clear:both;"></div></div></div><div class="module "><div class="modcontent clearfix"><p><a href="/oferta-academica/1769-nuevas-carreras"><img src="/images/NUEVASCARRERASok.jpg" alt="NUEVASCARRERASok.jpg" style="display: block; margin-left: auto; margin-right: auto;" /></a>&nbsp;</p><p><a href="/contenidoslideshow/53-proyecto-yo-me-sumo/2057-proyecto-transparencia"><img src="/images/YomeSumook.jpg" alt="YomeSumook.jpg" style="display: block; margin-left: auto; margin-right: auto;" /></a> <br /><br /></p></div></div></div></div></div></div></section><section id="yt_spotlight" class="block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="position-2" class="span12"><div class="module "><div class="modcontent clearfix"><div class="jmnewspro css3  layout9" id="jmnewspro-151"><div class="slider jm-bxslider" data-resize="1" data-useCSS="" data-mode="horizontal" data-easing="swing" data-slideSelector="" data-slideWidth="150" data-minSlides="1" data-maxSlides="20" data-moveSlides="0" data-slideMargin="10" data-autoHover="true" data-speed="500" data-adaptiveHeight="true" data-infiniteLoop="true" data-auto="false" data-pause="4000" data-controls="true" data-touchEnabled="1" data-onSliderLoad="jmnewspro151()" data-nextSelector="#jmnewspro-151 .jmnewspro-next" data-prevSelector="#jmnewspro-151 .jmnewspro-prev" data-nextText="Next" data-prevText="Prev"><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/989-educacion-virtual"><img src="/images/Educacion_Virtual218.jpg" alt="Educación Virtual"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/989-educacion-virtual">Educación Virtual</a></div><div class="slide-item-desc">Mat&iacute;as Virtual: Es el sistema de gesti&oacute;n de aprendizaje, la cual es utilizada para gestionar cursos en l&iacute;nea, as&iacute; como ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/989-educacion-virtual">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item image" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/663-evaluacion-docente"><img src="/images/Evaluac_Docente18.jpg" alt="Evaluación Docente "></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/663-evaluacion-docente">Evaluación Docente </a></div><div class="slide-item-desc">Estimado estudiante te notificamos que ya puedes completar la "Evaluaci&oacute;n Docente", tu participaci&oacute;n es clave para mejorar la docencia, ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/663-evaluacion-docente">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/188-conscius"><img src="/images/Conscius218.jpg" alt="Conscius"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/188-conscius">Conscius</a></div><div class="slide-item-desc">Conscius2: Es la nueva versi&oacute;n del sistema de gesti&oacute;n de aprendizaje institucional, la cual es utilizada para gestionar cursos en ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/188-conscius">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/189-uvirtual"><img src="/images/Uvirtual218.jpg" alt="Uvirtual"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/189-uvirtual">Uvirtual</a></div><div class="slide-item-desc">&nbsp;Puedes consultar: &nbsp;&gt; Calificaciones de tus materias inscritas &nbsp;&gt; Horarios de clases &nbsp;&gt; Evaluaci&oacute;n de tus ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/189-uvirtual">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/190-carreras-universitarias"><img src="/images/Careras_Universitarias18.jpg" alt="Carreras Universitarias"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/190-carreras-universitarias">Carreras Universitarias</a></div><div class="slide-item-desc">Te compartimos nuestra oferta acad&eacute;mica en carreras de pregrado, solo debes dar clic sobre el nombre de la carrera que deseas obtener ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/190-carreras-universitarias">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item image" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/ciclo-académico/horarios-de-clases"><img src="/images/Horarios_de_clases18.jpg" alt="Horarios de Clases"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/ciclo-académico/horarios-de-clases">Horarios de Clases</a></div><div class="slide-item-desc"> &nbsp; &nbsp; &nbsp; Te compartimos los horarios de clases, las cuales est&aacute;n clasificadas por Facultades y Escuelas.&nbsp;Solo debes ...</div> <span class="slide-item-readmore"><a target="_parent" href="/ciclo-académico/horarios-de-clases">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/ciclo-académico/cursos-de-formación-complementaria"><img src="/images/Cursos_Formac_Complementaria18.jpg" alt="Cursos de Formación Complementaria"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/ciclo-académico/cursos-de-formación-complementaria">Cursos de Formación Complementaria</a></div><div class="slide-item-desc"> Son requisito de graduaci&oacute;n y debes completarlos en el transcurso de tu carrera. Se imparten el transcurso de tu carrera. Se imparten ...</div> <span class="slide-item-readmore"><a target="_parent" href="/ciclo-académico/cursos-de-formación-complementaria">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/192-bolsa-de-trabajo-ujmd"><img src="/images/Bolsa_de_trabajo218.jpg" alt="Bolsa de Trabajo UJMD"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/192-bolsa-de-trabajo-ujmd">Bolsa de Trabajo UJMD</a></div><div class="slide-item-desc">La Bolsa de Trabajo de la Universidad Dr. Jos&eacute; Mat&iacute;as Delgado naci&oacute; con la misi&oacute;n de proveer un espacio de ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/192-bolsa-de-trabajo-ujmd">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/191-posgrados"><img src="/images/Posgrados_y_Educ_Continua18.jpg" alt="Posgrados y Educación Continua"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/191-posgrados">Posgrados y Educación Continua</a></div><div class="slide-item-desc">&gt;&nbsp;Conoce m&aacute;s aqu&iacute;</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/191-posgrados">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item image" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/ciclo-académico/horarios-de-inscripción"><img src="/images/Horarios_de_inscripcion218.jpg" alt="Horarios de Inscripción "></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/ciclo-académico/horarios-de-inscripción">Horarios de Inscripción </a></div><div class="slide-item-desc"> Te compartimos los horarios de inscripci&oacute;n en sus diferentes modalidades: &gt; En l&iacute;nea &gt; Presencial Solo debes dar clic en ...</div> <span class="slide-item-readmore"><a target="_parent" href="/ciclo-académico/horarios-de-inscripción">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/servicios-universitarios/servicios-de-la-universidad/informativo/catalogo-academico"><img src="/images/Catalogo_Estudiantil18.jpg" alt="Catálogo Académico "></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/servicios-universitarios/servicios-de-la-universidad/informativo/catalogo-academico">Catálogo Académico </a></div><div class="slide-item-desc">&nbsp;</div> <span class="slide-item-readmore"><a target="_parent" href="/servicios-universitarios/servicios-de-la-universidad/informativo/catalogo-academico">Leer más...</a></span> </div></div></div></div></div></div><div class="slide-item text" style="min-height:100px"><div class="slide-item-wrap"><div class="view slide-item-wrap-item"><div class="slide-item-image clearfix"> <a target="_parent" href="/banner-de-opciones/1239-juego-interactivo-papel-picado"><img src="/images/Papel_Picado18.jpg" alt="Juego Interactivo Papel Picado"></a> </div><div class="slide-item-desc-warp jmnewsprohover"><div class="slide-inner"><div class="padding"><div class="slide-item-title"><a target="_parent" href="/banner-de-opciones/1239-juego-interactivo-papel-picado">Juego Interactivo Papel Picado</a></div><div class="slide-item-desc"> Este juego es una aplicaci&oacute;n derivada del libro Un mundo en papel picado: Don Manuel Pasasin un Izalque&ntilde;o y su obra desarrollado por ...</div> <span class="slide-item-readmore"><a target="_parent" href="/banner-de-opciones/1239-juego-interactivo-papel-picado">Leer más...</a></span> </div></div></div></div></div></div></div><div class="NavButtons BottomRight clearfix"><div class="Inner"> <span class="jmnewspro-prev"></span> <span class="jmnewspro-next"></span> </div></div></div> <script type="text/javascript">function jmnewspro151(){}</script> </div> </div> </div> </div> </div> </div> </section><section id="content" class="content layout-mr block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="content_main" class="span9" data-normal="span9" data-tablet="span9" data-stablet="span9"><div class="content-main-inner "><div id="breadcrumb" class="span12" data-normal="span12" data-stablet="span12"><div class="module "><div class="modcontent clearfix"><table border="0" style="width: 728px;" align="center"> <tbody> <tr> <td style="width: 175px;"><img src="/images/Fotos_para_Contenido/bannerbibliteca.jpg" alt="bannerbibliteca" width="182" height="110" style="float: left;" /></td> <td>&nbsp;</td> <td style="width: 175px;"><img src="/images/Fotos_para_Contenido/REVISTAS.jpg" alt="REVISTAS" width="214" height="110" style="float: left;" /></td> <td>&nbsp;</td> <td><img src="/images/Fotos_para_Contenido/ASESORIA.jpg" alt="ASESORIA" width="165" height="110" style="float: left;" /></td> </tr> <tr> <td style="width: 175px;"><p><span style="color: #000080;"><strong><span style="font-family: arial, helvetica, sans-serif; font-size: 12pt;">BIBLIOTECA</span></strong></span></p><p><span style="font-family: arial, helvetica, sans-serif; font-size: 10pt;">La Biblioteca Universitaria Hugo Lindo, te ofrece los siguientes recursos: Bolet&iacute;n biblioteca, Sugerencias por especialidad, Documentos descargables, Herramientas de apoyo, e-recursos, etc.</span></p><p><a href="http://biblioteca.ujmd.edu.sv" target="_blank" style="font-family: arial, helvetica, sans-serif; font-size: 12pt;">Ingresar</a></p></td> <td>&nbsp;</td> <td style="width: 175px;" valign="top"><span style="color: #000080; font-size: 12pt;"><strong><span style="font-family: arial, helvetica, sans-serif;">REVISTAS DIGITALES</span></strong></span> <p>&nbsp;</p><p><span style="font-family: arial, helvetica, sans-serif; font-size: 10pt;">Ac&aacute; encontraras boletines especializados creados por las diferentes unidades acad&eacute;micas.</span></p><p>&nbsp;&nbsp;</p><p><a href="/investigación/revistas-digitales" style="font-family: arial, helvetica, sans-serif; font-size: 12pt;">Ingresar</a></p></td> <td>&nbsp;</td> <td style="width: 225px;" valign="top"><p><span style="color: #000080;"><strong><span style="font-family: arial, helvetica, sans-serif; font-size: 12pt;">Orientaci&oacute;n y Servicio al estudiante</span></strong></span></p><p><span style="font-family: arial, helvetica, sans-serif; font-size: 10pt;">La Universidad Dr. Jos&eacute; Mat&iacute;as Delgado en su af&aacute;n de prestar un mejor servicio a estudiantes activos y de nuevo ingreso, pone a tu disposici&oacute;n el servicio de Orientaci&oacute;n Vocacional y Educativa.</span></p><p>&nbsp;<a href="/index.php/la-universidad/unidades-de-apoyo-acad%C3%A9mico-administrativas/direcci%C3%B3n-de-orientaci%C3%B3n-y-servicio-al-estudiante" style="font-family: arial, helvetica, sans-serif; font-size: 12pt;">Leer m&aacute;s</a></p></td> </tr> </tbody> </table> </div> </div> </div><div class="span12 no-minheight"><div id="system-message-container"> </div> </div><div id="yt_component" class="span12" data-normal="" data-stablet=""><div class="component-inner"><div class="blog-featured"> </div> </div> </div><div id="position-5" class="span12" data-normal="span12" data-stablet="span12"><div class="module "><div class="modcontent clearfix"> ﻿ <script type="text/javascript">jQuery.noConflict();jQuery(function(){jQuery(document).ready(function()
{jQuery.noConflict();jQuery(function(){jQuery("#likebox_1").hover(function(){jQuery(this).stop(true,false).animate({right:0},500);},function(){jQuery("#likebox_1").stop(true,false).animate({right:-310},500);});jQuery("#polecam_1").hover(function(){jQuery(this).stop(true,false).animate({right:0},500);},function(){jQuery("#polecam_1").stop(true,false).animate({right:-310},500);});});});});</script><div id="likebox_1" style="right:-310px;top: 100px;"/><div id="likebox_1_1" style="text-align:left;width:300px;height:600px;"/><a class="open" id="fblink" href="#"></a><img style="margin-top: 25px;left:-38px;" src="/modules/mod_facebook_slide_likebox/tmpl/images/fb1.png" alt="" /><iframe src="http://www.facebook.com/plugins/likebox.php?id=117892388223741&amp;locale=es_LA&amp;width=300&amp;height=600&amp;colorscheme=light&amp;show_faces=true&amp;border_color&amp;stream=true&amp;header=false" scrolling="no" frameborder="0" style="border:none; overflow:hidden; width:300px; height:600px;" allowTransparency="true"></iframe></div></div><div id="polecam_1" style="top:100px; right:-310px;height:600px;"/><div id="polecam_1_1" style="width:300px;"/><a class="open" id="twlink" href="#"></a><img style="margin-top: 135px; left:-38px;" id="polecamy_img" src="/modules/mod_facebook_slide_likebox/tmpl/images/tw1.png"> <a class="twitter-timeline" width="300" height="600" data-theme="light" href="https://twitter.com/UJMD_sv" data-widget-id="348116677248049152">Tweets by @UJMD_sv</a> <script>!function(d,s,id){var js,fjs=d.getElementsByTagName(s)[0],p=/^http:/.test(d.location)?'http':'https';if(!d.getElementById(id)){js=d.createElement(s);js.id=id;js.src=p+"://platform.twitter.com/widgets.js";fjs.parentNode.insertBefore(js,fjs);}}(document,"script","twitter-wjs");</script> </div></div></div></div></div></div></div><div id="content_right" class="span3" data-normal="span3" data-tablet="span3" data-stablet="span3"><div class="content-right-in"><div id="position-7" class="span12" data-normal="" data-tablet="" data-stablet=""><div class="module "><h3 class="modtitle">Eventos </h3><div class="modcontent clearfix"><p><iframe src="https://www.facebook.com/plugins/page.php?href=https%3A%2F%2Fwww.facebook.com%2FUniversidadDrJoseMatiasDelgado%2F&amp;tabs=events&amp;width=320&amp;height=420&amp;small_header=true&amp;adapt_container_width=true&amp;hide_cover=true&amp;show_facepile=true&amp;appId" width="320" height="420" style="border: none; overflow: hidden; display: block; margin-left: auto; margin-right: auto;" frameborder="0" scrolling="no"></iframe></p></div></div><div class="module "><div class="modcontent clearfix"><p><a href="/la-universidad/todas-las-noticias"><img src="/images/Captura2.JPG" alt="Captura2" width="226" height="37" /></a></p></div></div></div></div></div></div></div></div></section><footer id="yt_footer" class="block"><div class="yt-main"><div class="yt-main-in1 container"><div class="yt-main-in2 row-fluid"><div id="yt_copyrightposition" class="span12"><div class="footer1">Copyright &#169; 2018 Universidad Dr. José Matías Delgado | El Salvador. All Rights Reserved. Designed by <a target="_blank" title="Visit SmartAddons!" href="http://www.smartaddons.com/">SmartAddons.Com</a></div><div class="footer2"></a> Campus 1: Km. 8 1/2 carretera a Santa Tecla. Tel. 2278-1011 o 2212-9400 Fax: 2289-5314 Campus 2: Calle el Pedregal y Av. Finca al Espino, frente a la entrada de Escuela Militar, Antiguo Cuscatlán. La Libertad.Facultad de Jurisprudencia y Ciencias Sociales Tel: 2241-7700. Fax 2289-4229 Facultad de Economía: Tel. 2212-9400 Fax. 2289-5314 Contáctenos:webmaster@ujmd.edu.sv </a></div></div></div></div></div></footer> <script type="text/javascript">jQuery(document).ready(function($){var headerbgimage='';var footerbgimage='';if(headerbgimage){$('#yt_header').addClass(headerbgimage);}});</script> <a id="yt-totop" class="backtotop" href="#"><i class="icon-chevron-up"></i></a> <script type="text/javascript">jQuery(".backtotop").addClass("hidden-top");jQuery(window).scroll(function(){if(jQuery(this).scrollTop()===0){jQuery(".backtotop").addClass("hidden-top")}else{jQuery(".backtotop").removeClass("hidden-top")}});jQuery('.backtotop').click(function(){jQuery('body,html').animate({scrollTop:0},1200);return false;});</script> </section> </body> </html>