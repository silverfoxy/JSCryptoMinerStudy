<!DOCTYPE html>
<!--[if lt IE 7 ]><html class="ie ie6" lang="es-ES"> <![endif]-->
<!--[if IE 7 ]><html class="ie ie7" lang="es-ES"> <![endif]-->
<!--[if IE 8 ]><html class="ie ie8" lang="es-ES"> <![endif]-->
<!--[if IE 9 ]><html class="ie ie9" lang="es-ES"> <![endif]-->
<!--[if !(IE)]><!--><html lang="es-ES"> <!--<![endif]-->
<head><link rel="stylesheet" type="text/css" href="http://ultimahora.sv/wp-content/cache/minify/7091a.css" media="all" />

      <!-- Basic Page Needs
  	  ================================================== -->
	<meta charset="UTF-8" />
	<meta http-equiv="content-type" content="text/html; charset=UTF-8">
	<meta name="google-site-verification" content="ZQJtqEXDtnLNfUq7NMh4SoV3UoObJSgKDNlNxYG2AZ4" />
    <meta property="fb:pages" content="1524382234487630">
    <title>Última Hora SV | Un periódico con información para los que no se detienen</title>
        <!-- Mobile Specific Metas
  		================================================== -->
           <meta name="viewport" content="width=device-width, initial-scale=1.0">
        <!-- Favicons
        ================================================== -->
                    <link rel="shortcut icon" href="http://ultimahora.sv/wp-content/uploads/2016/10/faviconuh.png" type="image/x-icon" />       
    
<title>Última Hora SV</title>

<!-- Inicio The SEO Framework por Sybre Waaijer -->
<meta name="robots" content="noydir" />
<meta name="description" content="Un periódico con información para los que no se detienen en" />
<meta property="og:image" content="" />
<meta property="og:locale" content="es_ES" />
<meta property="og:type" content="website" />
<meta property="og:title" content="Última Hora SV" />
<meta property="og:description" content="Un periódico con información para los que no se detienen en" />
<meta property="og:url" content="http://ultimahora.sv/" />
<link rel="canonical" href="http://ultimahora.sv/" />
<script type="application/ld+json">{"@context":"http://schema.org","@type":"WebSite","url":"http://ultimahora.sv/","potentialAction":{"@type":"SearchAction","target":"http://ultimahora.sv/search/{search_term_string}","query-input":"required name=search_term_string"}}</script>
<script type="application/ld+json">{"@context":"http://schema.org","@type":"Organization","url":"http://ultimahora.sv/"}</script>
<!-- Final The SEO Framework por Sybre Waaijer | 0.00011s -->

<link rel='dns-prefetch' href='//platform.twitter.com' />
<link rel='dns-prefetch' href='//fonts.googleapis.com' />
<link rel='dns-prefetch' href='//s.w.org' />
<link rel="alternate" type="application/rss+xml" title=" &raquo; Feed" href="http://ultimahora.sv/feed/" />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.3\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.3\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/ultimahora.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.8.5"}};
			!function(a,b,c){function d(a){var b,c,d,e,f=String.fromCharCode;if(!k||!k.fillText)return!1;switch(k.clearRect(0,0,j.width,j.height),k.textBaseline="top",k.font="600 32px Arial",a){case"flag":return k.fillText(f(55356,56826,55356,56819),0,0),b=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,56826,8203,55356,56819),0,0),c=j.toDataURL(),b!==c&&(k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57332,56128,56423,56128,56418,56128,56421,56128,56430,56128,56423,56128,56447),0,0),b=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57332,8203,56128,56423,8203,56128,56418,8203,56128,56421,8203,56128,56430,8203,56128,56423,8203,56128,56447),0,0),c=j.toDataURL(),b!==c);case"emoji4":return k.fillText(f(55358,56794,8205,9794,65039),0,0),d=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55358,56794,8203,9794,65039),0,0),e=j.toDataURL(),d!==e}return!1}function e(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var f,g,h,i,j=b.createElement("canvas"),k=j.getContext&&j.getContext("2d");for(i=Array("flag","emoji4"),c.supports={everything:!0,everythingExceptFlag:!0},h=0;h<i.length;h++)c.supports[i[h]]=d(i[h]),c.supports.everything=c.supports.everything&&c.supports[i[h]],"flag"!==i[h]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[i[h]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(g=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",g,!1),a.addEventListener("load",g,!1)):(a.attachEvent("onload",g),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),f=c.source||{},f.concatemoji?e(f.concatemoji):f.wpemoji&&f.twemoji&&(e(f.twemoji),e(f.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>









<link rel='stylesheet' id='nanomag_fonts_url-css'  href='//fonts.googleapis.com/css?family=Open+Sans%3A300%2C400%2C600%2C700%2C800%2C900%2C400italic%2C700italic%2C900italic%7COpen+Sans%3A300%2C400%2C600%2C700%2C800%2C900%2C400italic%2C700italic%2C900italic%7COpen+Sans%3A300%2C400%2C600%2C700%2C800%2C900%2C400italic%2C700italic%2C900italic%7COpen+Sans%3A300%2C400%2C600%2C700%2C800%2C900%2C400italic%2C700italic%2C900italic%7C&#038;subset=latin%2Clatin-ext%2Ccyrillic%2Ccyrillic-ext%2Cgreek%2Cgreek-ext%2Cvietnamese&#038;ver=1.0.0' type='text/css' media='all' />







<link rel='stylesheet' id='nanomag_custom-style-css'  href='http://ultimahora.sv/wp-content/themes/nanomag/custom_style.php?ver=1.6' type='text/css' media='all' />

<style id='__EPYT__style-inline-css' type='text/css'>

                .epyt-gallery-thumb {
                        width: 33.333%;
                }
                
</style>
<script type='text/javascript'>
/* <![CDATA[ */
var user_review_script = {"post_id":"5","ajaxurl":"http:\/\/ultimahora.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/b2fe6.js"></script>



<script type='text/javascript'>
/* <![CDATA[ */
var bwg_objectsL10n = {"bwg_select_tag":"Select Tag","bwg_search":"Buscar"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/f8880.js"></script>




<script type='text/javascript'>
/* <![CDATA[ */
var bwg_objectL10n = {"bwg_field_required":"se requiere el campo. ","bwg_mail_validation":"Esta no es una direcci\u00f3n de correo electr\u00f3nico v\u00e1lida.","bwg_search_result":"No hay im\u00e1genes que coincidan con su b\u00fasqueda."};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/4a079.js"></script>


<script type='text/javascript'>
/* <![CDATA[ */
var _EPYT_ = {"ajaxurl":"http:\/\/ultimahora.sv\/wp-admin\/admin-ajax.php","security":"fe2275fa76","gallery_scrolloffset":"20","eppathtoscripts":"http:\/\/ultimahora.sv\/wp-content\/plugins\/youtube-embed-plus\/scripts\/","epresponsiveselector":"[\"iframe.__youtube_prefs_widget__\"]","epdovol":"1","version":"11.8.6.1","evselector":"iframe.__youtube_prefs__[src], iframe[src*=\"youtube.com\/embed\/\"], iframe[src*=\"youtube-nocookie.com\/embed\/\"]","ajax_compat":"","stopMobileBuffer":"1"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/8fc7a.js"></script>

<link rel='https://api.w.org/' href='http://ultimahora.sv/wp-json/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://ultimahora.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://ultimahora.sv/wp-includes/wlwmanifest.xml" /> 
<link rel="alternate" type="application/json+oembed" href="http://ultimahora.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fultimahora.sv%2F" />
<link rel="alternate" type="text/xml+oembed" href="http://ultimahora.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fultimahora.sv%2F&#038;format=xml" />

<!-- This site is using AdRotate v4.10 to display their advertisements - https://ajdg.solutions/products/adrotate-for-wordpress/ -->
<!-- afb Instant Articles -->
			<meta property="fb:pages" content="1524382234487630" /><meta property="fb:app_id" content="271202853384837"/><!--[if lt IE 9]><script src="http://html5shim.googlecode.com/svn/trunk/html5.js"></script><![endif]-->
    <meta name="twitter:widgets:link-color" content="#000000" /><meta name="twitter:widgets:border-color" content="#000000" /><meta name="twitter:partner" content="tfwp" />
<meta name="twitter:card" content="summary" /><meta name="twitter:site" content="@ultimahsv" /><meta name="twitter:description" content="Un periódico con información para los que no se detienen" />
<script async src="//pagead2.googlesyndication.com/pagead/js/adsbygoogle.js"></script>
<script>
  (adsbygoogle = window.adsbygoogle || []).push({
    google_ad_client: "ca-pub-2104763040190014",
    enable_page_level_ads: true
  });
</script>
<!-- end head -->
</head>
<body class="home page-template page-template-home-page page-template-home-page-php page page-id-5 magazine_default_layout" itemscope="itemscope" itemtype="http://schema.org/WebPage">
   
<div id="sb-site" class="body_wraper_full">     			

        <!-- Start header -->

<!-- Header6 layout --> 

<header class="header-wraper theme_header_style_5">

<div class="header_top_wrapper">
<div class="row">
<div class="six columns header-top-left-bar">

              <div class="news_ticker_wrapper">
<div class="row">
<div class="twelve columns">
  <div id="ticker">
  <div class="tickerfloat_wrapper"><div class="tickerfloat">Noticias de Última Hora</div></div>
   <div class="marquee" id="mycrawler">
           
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/">Jaime “La Chelona” Rodríguez acusado de malversación de fondos</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/">GANA presenta a la Fiscalía aviso de fraude electoral en San Vicente</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/">Alcaldía de Santa Tecla instala 6 cámaras de videovigilancia en bulevar Monseñor Romero</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/fiscalia-insiste-en-quitarle-patrimonio-familiar-a-diputado-cardoza/">Fiscalía insiste en quitarle patrimonio familiar a diputado Cardoza</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/">Jefe de Sección de Probidad busca formar parte de Sala de lo Constitucional</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/renuncia-presidente-de-peru/">Renuncia presidente de Perú</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/reynaldo-cardoza-aspira-una-vicepresidencia-o-la-presidencia-de-asamblea/">Reynaldo Cardoza aspira una vicepresidencia o la presidencia de Asamblea</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/partidos-politicos-inician-cabildeo-por-presidencia-de-asamblea-legislativa/">Partidos políticos inician cabildeo por presidencia de Asamblea Legislativa</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/ortiz-renuncia-a-sus-aspiraciones-presidenciales/">Ortiz renuncia a sus aspiraciones presidenciales</a>
      </div>

            
       <div>
        <span class="ticker_dot"><i class="fa fa-chevron-right"></i></span><a class="ticker_title" href="http://ultimahora.sv/interiano-asegura-que-arena-logro-una-gran-campana-con-bajo-presupuesto/">Interiano asegura que ARENA logró una gran campaña con bajo presupuesto</a>
      </div>

                
        </div>
        </div>
    
</div>

</div>
</div>
    
</div>

<div class="six columns header-top-right-bar">

<a class="open toggle-lef sb-toggle-left navbar-left" href="#nav">
        <div class="navicon-line"></div>
        <div class="navicon-line"></div>
        <div class="navicon-line"></div>
        </a>
      <div id="search_block_top">
    <form id="searchbox" action="http://ultimahora.sv/" method="GET" role="search">
        <p>
            <input type="text" id="search_query_top" name="s" class="search_query ac_input" value="" placeholder="Buscar">
           <button type="submit"><i class="fa fa-search"></i></button>
    </p>
    </form>
    <span>Search</span>
    <div class="clearfix"></div>
</div>


  
    <ul class="social-icons-list top-bar-social">
      <li><a href="https://www.facebook.com/ultimahsv" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/facebook.png" alt="Facebook"></a></li>                    <li><a href="https://www.youtube.com/channel/UCxD1dNdPTM7LxkghZ_5wFrA" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/youtube.png" alt="Youtube"></a></li>                    <li><a href="https://twitter.com/ultimahsv" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/twitter.png" alt="Twitter"></a></li>                                                     </ul>  
      
<div class="clearfix"></div>
</div>

</div>
</div>

 
        
 <div class="header_main_wrapper"> 
        <div class="row">
    <div class="four columns header-top-left">
    
      <!-- begin logo -->
                           
                           
                                <a href="http://ultimahora.sv/">
                                                                           
                                        <img src="http://ultimahora.sv/wp-content/uploads/2016/09/logofront.png" alt="Un periódico con información para los que no se detienen" id="theme_logo_img" />
                                                                    </a>
                            
                            <!-- end logo -->
    </div>
        <div class="eight columns header-top-right">  
  <div class="textwidget custom-html-widget"><div class="centered" style="width: 100%;height: 90%;text-align: center;m;margin-top: 15px;">   
    <a href="http://ultimahora.sv/category/arena/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/ARENA-1.png" style="width: 10%;height: auto;margin-right: 10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/fmln/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/FMLN-1.png" style="width: 10%;height: auto;margin-right: 10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/gana/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/GANA-1.jpg" style="width: 10%;height: auto;margin-right: 10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/pcn/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/PCN-1.jpg" style="width: 10%;height: auto;margin-right: 10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/pdc/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/PDC-1.jpg" style="width: 10%;height: auto;margin-right:10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/cd/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/08/CD.jpg" style="width: 10%;height: auto;margin-right:10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/nuevas-ideas/">
        <img src="http://ultimahora.sv/wp-content/uploads/2018/01/nuevas_ideas.png" style="width: 10%;height: auto;margin-right:10px;/* border-radius: 5px; */">
    </a>
    <a href="http://ultimahora.sv/category/clase-politica/encuestas/">
        <img src="http://ultimahora.sv/wp-content/uploads/2017/09/BOTON.jpg" style="width: 10%;height: auto; /* border-radius: 5px; */">
    </a>
</div></div>    </div>
        
</div>

</div>

                
<!-- end header, logo, top ads -->

              
<!-- Start Main menu -->
<div id="menu_wrapper" class="menu_wrapper ">
<div class="menu_border_top_full"></div>
<div class="row">
    <div class="main_menu twelve columns"> 
        <div class="menu_border_top"></div>
                            <!-- main menu -->
                           
  <div class="menu-primary-container main-menu">
<ul id="mainmenu" class="sf-menu"><li id="menu-item-17" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children"><a href="http://ultimahora.sv/category/portada/portada-portada/">portada<span class="border-menu"></span></a><ul class="sub-menu">	<li id="menu-item-20" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/portada/portada-portada/politica/">Política<span class="border-menu"></span></a></li>

					</ul></li>
<li id="menu-item-14" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/economia/">Economía<span class="border-menu"></span></a></li>
<li id="menu-item-7913" class="menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/negocios/">Negocios<span class="border-menu"></span></a></li>
<li id="menu-item-16" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children"><a href="http://ultimahora.sv/category/internacionales/">Internacionales<span class="border-menu"></span></a><ul class="sub-menu">	<li id="menu-item-25" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento<span class="border-menu"></span></a></li>
	<li id="menu-item-22" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/internacionales/tecnologia/">Tecnología<span class="border-menu"></span></a></li>

					</ul></li>
<li id="menu-item-24" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/internacionales/deportes/">Deportes<span class="border-menu"></span></a></li>
<li id="menu-item-13" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children"><a href="http://ultimahora.sv/category/clase-politica/">Clase política<span class="border-menu"></span></a><ul class="sub-menu">	<li id="menu-item-15" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/editoriales/">Editoriales<span class="border-menu"></span></a></li>
	<li id="menu-item-23" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/editoriales/especiales/">Especiales<span class="border-menu"></span></a></li>
	<li id="menu-item-26" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/clase-politica/encuestas/">Encuestas<span class="border-menu"></span></a></li>

					</ul></li>
<li id="menu-item-18" class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana<span class="border-menu"></span></a></li>
<li id="menu-item-66763" class="menu-item menu-item-type-post_type menu-item-object-page"><a href="http://ultimahora.sv/tv/">UH TV<span class="border-menu"></span></a></li>
</ul><div class="clearfix"></div>
</div>                             
                            <!-- end main menu -->                                                                                   
                        </div>                                           
                    </div>   
                    </div>
            </header>



  
<div id="content_nav">
        <div id="nav">
        <ul id="mobile_menu_slide" class="menu_moble_slide"><li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children menu-item-17"><a href="http://ultimahora.sv/category/portada/portada-portada/">portada<span class="border-menu"></span></a>
<ul  class="sub-menu">
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-20"><a href="http://ultimahora.sv/category/portada/portada-portada/politica/">Política<span class="border-menu"></span></a></li>
</ul>
</li>
<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-14"><a href="http://ultimahora.sv/category/economia/">Economía<span class="border-menu"></span></a></li>
<li class="menu-item menu-item-type-taxonomy menu-item-object-category menu-item-7913"><a href="http://ultimahora.sv/category/negocios/">Negocios<span class="border-menu"></span></a></li>
<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children menu-item-16"><a href="http://ultimahora.sv/category/internacionales/">Internacionales<span class="border-menu"></span></a>
<ul  class="sub-menu">
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-25"><a href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento<span class="border-menu"></span></a></li>
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-22"><a href="http://ultimahora.sv/category/internacionales/tecnologia/">Tecnología<span class="border-menu"></span></a></li>
</ul>
</li>
<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-24"><a href="http://ultimahora.sv/category/internacionales/deportes/">Deportes<span class="border-menu"></span></a></li>
<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-has-children menu-item-13"><a href="http://ultimahora.sv/category/clase-politica/">Clase política<span class="border-menu"></span></a>
<ul  class="sub-menu">
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-15"><a href="http://ultimahora.sv/category/editoriales/">Editoriales<span class="border-menu"></span></a></li>
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-23"><a href="http://ultimahora.sv/category/editoriales/especiales/">Especiales<span class="border-menu"></span></a></li>
	<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-26"><a href="http://ultimahora.sv/category/clase-politica/encuestas/">Encuestas<span class="border-menu"></span></a></li>
</ul>
</li>
<li class="megamenu columns-3 color-2 menu-item menu-item-type-taxonomy menu-item-object-category menu-item-18"><a href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana<span class="border-menu"></span></a></li>
<li class="menu-item menu-item-type-post_type menu-item-object-page menu-item-66763"><a href="http://ultimahora.sv/tv/">UH TV<span class="border-menu"></span></a></li>
</ul>   </div>
    </div>             
<div class="slider_wrapper_main">
<div class="row header-slider-home header-slider-home-list-right">
  <div class="twelve columns feature-three"> 
  <div class="slide-large-wrapper header-slider2">
      <div class="owl_slider slider-large owl-carousel">
            
 
<div class="item_slide">
<div class="main-post-image-slider image_post">
<a href="http://ultimahora.sv/ortiz-renuncia-a-sus-aspiraciones-presidenciales/" class="feature-link" title="Ortiz renuncia a sus aspiraciones presidenciales">              
<img width="640" height="399" src="http://ultimahora.sv/wp-content/uploads/2018/03/oscar-ortiz.jpg" class="attachment-slider-normal size-slider-normal wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/oscar-ortiz.jpg 640w, http://ultimahora.sv/wp-content/uploads/2018/03/oscar-ortiz-300x187.jpg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/oscar-ortiz-171x108.jpg 171w" sizes="(max-width: 640px) 100vw, 640px" /> 
</a>
<div class="item_slide_caption">
 <p class="post-meta meta-main-img"><span class="post-date updated"><i class="fa fa-clock-o"></i>Mar 21, 2018</span><span class="meta-cat"><i class="fa fa-folder-o"></i><a href="http://ultimahora.sv/category/clase-politica/" rel="category tag">Clase política</a>, <a href="http://ultimahora.sv/category/fmln/" rel="category tag">FMLN</a>, <a href="http://ultimahora.sv/category/portada/" rel="category tag">Portada</a></span></p>                                <h1><a class="heading" href="http://ultimahora.sv/ortiz-renuncia-a-sus-aspiraciones-presidenciales/">Ortiz renuncia a sus aspiraciones presidenciales</a> </h1>                                              
            </div>
</div>
              
                      
<div class="sub-post-image-slider image_post">
<a href="http://ultimahora.sv/felix-ulloa-el-partido-nuevas-ideas-ya-existe/" class="feature-link" title="Félix Ulloa: El partido Nuevas Ideas ya existe">              
<img width="240" height="140" src="http://ultimahora.sv/wp-content/uploads/2018/03/DY0Fm5xX0AUqCUr-240x140.jpg" class="attachment-slider-small size-slider-small wp-post-image" alt="" /></a>

<div class="item_slide_caption">
                                <h1><a href="http://ultimahora.sv/felix-ulloa-el-partido-nuevas-ideas-ya-existe/">Félix Ulloa: El partido Nuevas Ideas ya existe</a> </h1>
                                                                                     
            </div>

</div>
              
                      
<div class="sub-post-image-slider image_post">
<a href="http://ultimahora.sv/hugo-martinez-los-partidos-deben-renovarse-para-no-poner-en-crisis-el-sistema-politico/" class="feature-link" title="Hugo Martínez: Los partidos deben renovarse para no poner en crisis el sistema político">              
<img width="240" height="140" src="http://ultimahora.sv/wp-content/uploads/2018/03/hugo-martinez-e1521638505476-240x140.jpg" class="attachment-slider-small size-slider-small wp-post-image" alt="" /></a>

<div class="item_slide_caption">
                                <h1><a href="http://ultimahora.sv/hugo-martinez-los-partidos-deben-renovarse-para-no-poner-en-crisis-el-sistema-politico/">Hugo Martínez: Los partidos deben renovarse para no poner en crisis el sistema político</a> </h1>
                                                                                     
            </div>

</div>
              
                      
<div class="sub-post-image-slider image_post">
<a href="http://ultimahora.sv/dagoberto-gutierrez-en-el-gobierno-hay-desesperacion-dispersion-y-decepcion/" class="feature-link" title="Dagoberto Gutiérrez: En el Gobierno hay desesperación, dispersión y decepción">              
<img width="240" height="140" src="http://ultimahora.sv/wp-content/uploads/2018/03/DYvK2YFVoAIC1MX-240x140.jpg" class="attachment-slider-small size-slider-small wp-post-image" alt="" /></a>

<div class="item_slide_caption">
                                <h1><a href="http://ultimahora.sv/dagoberto-gutierrez-en-el-gobierno-hay-desesperacion-dispersion-y-decepcion/">Dagoberto Gutiérrez: En el Gobierno hay desesperación, dispersión y decepción</a> </h1>
                                                                                     
            </div>

</div>
              
                             </div>  
               
                
                   
              </div>
 </div>
  <div class="slider-right-list-post">
<h2 class="right-list-post-title">Editoriales</h2>

                      <ul class="feature-post-list scroll_list_post">  
                    
<li>
<a  href="http://ultimahora.sv/goku-veni-en-nombre-de-el-salvador/" class="feature-image-link image_post" title="Gokú, vení en nombre de El Salvador">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/35c28593-ae25-4c14-8d21-81977533688e-100x75.jpeg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/goku-veni-en-nombre-de-el-salvador/">Gokú, vení en nombre de El Salvador</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 19, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/renuncie-senor-olivo/" class="feature-image-link image_post" title="Renuncie, señor Olivo">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/TSE-Partidos-28082014_16-770x438-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/renuncie-senor-olivo/">Renuncie, señor Olivo</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 18, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/uhtv-analisis-juan-valiente/" class="feature-image-link image_post" title="#UHTV | Análisis Juan Valiente">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Captura-de-pantalla-2018-03-15-a-las-10.17.04-100x75.png" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/uhtv-analisis-juan-valiente/">#UHTV | Análisis Juan Valiente</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 15, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/revolucion-o-muerte/" class="feature-image-link image_post" title="¡Revolución o Muerte!">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/d8689ef2-f76e-4ac6-97d8-fa9561a3faa5-100x75.jpeg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a><a class="post-category-color-text" style="color:#f34035" href="http://ultimahora.sv/category/portada/">Portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/revolucion-o-muerte/">¡Revolución o Muerte!</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 09, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/dios-y-la-politica/" class="feature-image-link image_post" title="Dios y la política">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/MG_6309-e1520119901996-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/dios-y-la-politica/">Dios y la política</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 03, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/un-candidato-que-no-quiere-debatir-es-porque-tiene-poco-que-proponer-y-mucho-que-esconder/" class="feature-image-link image_post" title="Un candidato que no quiere debatir es porque tiene poco que proponer y mucho que esconder">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/01/IMG-20180108-WA0000-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a><a class="post-category-color-text" style="color:#f34035" href="http://ultimahora.sv/category/portada/">Portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/un-candidato-que-no-quiere-debatir-es-porque-tiene-poco-que-proponer-y-mucho-que-esconder/">Un candidato que no quiere debatir es porque tiene poco que proponer y mucho que esconder</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 08, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

                
<li>
<a  href="http://ultimahora.sv/10-deseos-para-el-salvador-en-el-2018/" class="feature-image-link image_post" title="10 deseos para El Salvador en el 2018">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/12/Bandera-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
  <span class="meta-category-small"><a class="post-category-color-text" style="color:#81d742" href="http://ultimahora.sv/category/editoriales/">Editoriales</a><a class="post-category-color-text" style="color:#f34035" href="http://ultimahora.sv/category/portada/">Portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/10-deseos-para-el-salvador-en-el-2018/">10 deseos para El Salvador en el 2018</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 01, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>

       
        
      </ul>
            </div>  
    </div>
    </div>
  </div>


<div class="carousel_post_home_wrapper">
<div class="row carousel_post_home">
  <div class="twelve columns carousel_header_wrapper">
 <div class="widget-title"><h2>Lo último</h2></div>  
  
 <div class="owl_carousel carousel_header">
 
 
                
 <div class="item carousel_header_medium ">
  
  <div class="two-content-wrapper medium-two-columns ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/" class="feature-link" title="Jaime “La Chelona” Rodríguez acusado de malversación de fondos">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Rodríguez-1-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
 
 <h3 class="image-post-title"><a href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/">Jaime “La Chelona” Rodríguez acusado de malversación de fondos</a></h3>      
 <p class="car_header_desc">El Juzgado 9° de Instrucción recibió de la Fiscalía General de la República la... </p>
 <div class="footer_meta"><a href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

 </div>
          
 <div class="item carousel_header_medium ">
  
  <div class="two-content-wrapper medium-two-columns ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/" class="feature-link" title="GANA presenta a la Fiscalía aviso de fraude electoral en San Vicente">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/GANA-Fiscalía-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
 
 <h3 class="image-post-title"><a href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/">GANA presenta a la Fiscalía aviso de fraude electoral en San Vicente</a></h3>      
 <p class="car_header_desc">El diputado de GANA, Juan Pablo Herrera presentó un aviso por fraude electoral en el... </p>
 <div class="footer_meta"><a href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

 </div>
          
 <div class="item carousel_header_medium ">
  
  <div class="two-content-wrapper medium-two-columns ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/" class="feature-link" title="Jefe de Sección de Probidad busca formar parte de Sala de lo Constitucional">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/get_img-e1521666339866-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
 
 <h3 class="image-post-title"><a href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/">Jefe de Sección de Probidad busca formar parte de Sala de lo Constitucional</a></h3>      
 <p class="car_header_desc">El jefe de Sección de Probidad de la Corte Suprema de Justicia, Carlos Pineda busca una... </p>
 <div class="footer_meta"><a href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

 </div>
    

 
  </div>
  </div>
</div>
</div>


<!-- Start content -->
<div class="row main_content">
<div class="content_wraper three_columns_container">
   <!-- Start content -->
     <div class="eight columns content_display_col1" id="content">
            
			  <div id="aq-template-wrapper-44" class="aq-template-wrapper aq_row"><div id="aq-block-44-1" class="aq-block aq-block-home_large_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-8">
        <div class="widget-title"><h2>Nacionales</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="post_list_medium_widget"> 
    <div class="feature-post-list list-post-builder loop-post-content list-with-below-grid ">    
    <div class="image_post feature-item grid_below_image">
                 <a href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/" class="feature-link" title="Alcaldía de Santa Tecla instala 6 cámaras de videovigilancia en bulevar Monseñor Romero">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Alcaldia-Santa-Tecla-e1521673575951-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="post_loop_content">
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67318" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>    
 <h3 class="image-post-title feature_2col"><a href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/">Alcaldía de Santa Tecla instala 6 cámaras de videovigilancia en bulevar Monseñor Romero</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p><p class="post_des">El alcalde de Santa Tecla, Roberto d’Aubuisson, instaló seis nuevas cámaras de videovigilancia en el bulevar Monseñor Arnulfo Romero, esto como parte del proyecto... </p>
<a class="more_button_post" href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/">Leer más</a>
</div>
 </div>
    </div>



     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow">   
                					
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/fiscalia-insiste-en-quitarle-patrimonio-familiar-a-diputado-cardoza/" class="feature-image-link image_post" title="Fiscalía insiste en quitarle patrimonio familiar a diputado Cardoza">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/FGR-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/FGR-100x75.jpg 100w, http://ultimahora.sv/wp-content/uploads/2018/03/FGR-300x225.jpg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/FGR-768x576.jpg 768w, http://ultimahora.sv/wp-content/uploads/2018/03/FGR-1024x768.jpg 1024w, http://ultimahora.sv/wp-content/uploads/2018/03/FGR.jpg 1040w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/nacionales/">Nacionales</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/fiscalia-insiste-en-quitarle-patrimonio-familiar-a-diputado-cardoza/">Fiscalía insiste en quitarle patrimonio familiar a diputado Cardoza</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/representante-de-la-onu-pide-no-prorrogar-medidas-extraordinarias/" class="feature-image-link image_post" title="Representante de la ONU pide no prorrogar medidas extraordinarias">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/callamard-onu-pnc-sv-100x75.png" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/nacionales/">Nacionales</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/uncategorized/">Uncategorized</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/representante-de-la-onu-pide-no-prorrogar-medidas-extraordinarias/">Representante de la ONU pide no prorrogar medidas extraordinarias</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/medidas-extraordinarias-no-son-aprobadas-por-falta-de-consenso/" class="feature-image-link image_post" title="Medidas extraordinarias no son aprobadas por falta de consenso">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/plenaria-100x75.jpeg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/plenaria-100x75.jpeg 100w, http://ultimahora.sv/wp-content/uploads/2018/03/plenaria-300x225.jpeg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/plenaria-768x576.jpeg 768w, http://ultimahora.sv/wp-content/uploads/2018/03/plenaria-1024x768.jpeg 1024w, http://ultimahora.sv/wp-content/uploads/2018/03/plenaria.jpeg 1152w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/nacionales/">Nacionales</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/uncategorized/">Uncategorized</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/medidas-extraordinarias-no-son-aprobadas-por-falta-de-consenso/">Medidas extraordinarias no son aprobadas por falta de consenso</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/camara-especializada-ordena-repetir-el-juicio-del-caso-tregua-entre-pandillas/" class="feature-image-link image_post" title="Cámara especializada ordena repetir el juicio del caso tregua entre pandillas">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/05/caso-tregua-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/camara-especializada-ordena-repetir-el-juicio-del-caso-tregua-entre-pandillas/">Cámara especializada ordena repetir el juicio del caso tregua entre pandillas</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/presidente-sanchez-ceren-juramenta-a-nuevos-funcionarios/" class="feature-image-link image_post" title="Presidente Sánchez Cerén juramenta a nuevos funcionarios">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Juramenta-nuevos-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/presidente-sanchez-ceren-juramenta-a-nuevos-funcionarios/">Presidente Sánchez Cerén juramenta a nuevos funcionarios</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/alejandrina-castro-debe-trabajarse-por-un-estatus-migratorio-permanente/" class="feature-image-link image_post" title="Alejandrina Castro: Debe trabajarse por un estatus migratorio permanente">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Alejandrina-Castro-e1521491654327-100x75.jpeg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/nacionales/">Nacionales</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/alejandrina-castro-debe-trabajarse-por-un-estatus-migratorio-permanente/">Alejandrina Castro: Debe trabajarse por un estatus migratorio permanente</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 19, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-2" class="aq-block aq-block-aq_text_block aq_span12 aq-first clearfix"><p><a href="http://www.fedecredito.com.sv" target="_blank"><img src="http://ultimahora.sv/wp-content/uploads/2018/01/banner-fede.gif" class="img-responsive"></a></p>
</div><div id="aq-block-44-3" class="aq-block aq-block-home_large_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-8">
        <div class="widget-title"><h2>Clase política</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="post_list_medium_widget"> 
    <div class="feature-post-list list-post-builder loop-post-content list-with-below-grid ">    
    <div class="image_post feature-item grid_below_image">
                 <a href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/" class="feature-link" title="Jaime “La Chelona” Rodríguez acusado de malversación de fondos">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Rodríguez-1-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="post_loop_content">
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#ff3a3a" href="http://ultimahora.sv/category/fmln/">FMLN</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67326" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>    
 <h3 class="image-post-title feature_2col"><a href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/">Jaime “La Chelona” Rodríguez acusado de malversación de fondos</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p><p class="post_des">El Juzgado 9° de Instrucción recibió de la Fiscalía General de la República la acusación en contra de Jaime “La Chelona” Rodríguez por el delito de... </p>
<a class="more_button_post" href="http://ultimahora.sv/jaime-la-chelona-rodriguez-acusado-de-malversacion-de-fondos/">Leer más</a>
</div>
 </div>
    </div>



     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow">   
                					
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/" class="feature-image-link image_post" title="GANA presenta a la Fiscalía aviso de fraude electoral en San Vicente">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/GANA-Fiscalía-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#ff9000" href="http://ultimahora.sv/category/gana/">GANA</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/gana-presenta-a-la-fiscalia-aviso-de-fraude-electoral-en-san-vicente/">GANA presenta a la Fiscalía aviso de fraude electoral en San Vicente</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/" class="feature-image-link image_post" title="Jefe de Sección de Probidad busca formar parte de Sala de lo Constitucional">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/get_img-e1521666339866-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/jefe-de-seccion-de-probidad-busca-formar-parte-de-sala-de-lo-constitucional/">Jefe de Sección de Probidad busca formar parte de Sala de lo Constitucional</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/reynaldo-cardoza-aspira-una-vicepresidencia-o-la-presidencia-de-asamblea/" class="feature-image-link image_post" title="Reynaldo Cardoza aspira una vicepresidencia o la presidencia de Asamblea">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/02/REynaldo-Cardoza-e1519181971883-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/reynaldo-cardoza-aspira-una-vicepresidencia-o-la-presidencia-de-asamblea/">Reynaldo Cardoza aspira una vicepresidencia o la presidencia de Asamblea</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/partidos-politicos-inician-cabildeo-por-presidencia-de-asamblea-legislativa/" class="feature-image-link image_post" title="Partidos políticos inician cabildeo por presidencia de Asamblea Legislativa">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/02/Asamblea140220131-e1486647393404-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#ff9000" href="http://ultimahora.sv/category/gana/">GANA</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/partidos-politicos-inician-cabildeo-por-presidencia-de-asamblea-legislativa/">Partidos políticos inician cabildeo por presidencia de Asamblea Legislativa</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/ortiz-renuncia-a-sus-aspiraciones-presidenciales/" class="feature-image-link image_post" title="Ortiz renuncia a sus aspiraciones presidenciales">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/oscar-ortiz-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#ff3a3a" href="http://ultimahora.sv/category/fmln/">FMLN</a><a class="post-category-color-text" style="color:#f34035" href="http://ultimahora.sv/category/portada/">Portada</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/ortiz-renuncia-a-sus-aspiraciones-presidenciales/">Ortiz renuncia a sus aspiraciones presidenciales</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/interiano-asegura-que-arena-logro-una-gran-campana-con-bajo-presupuesto/" class="feature-image-link image_post" title="Interiano asegura que ARENA logró una gran campaña con bajo presupuesto">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/mauricio-interiano-e1521651748383-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/interiano-asegura-que-arena-logro-una-gran-campana-con-bajo-presupuesto/">Interiano asegura que ARENA logró una gran campaña con bajo presupuesto</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-4" class="aq-block aq-block-home_large_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-8">
        <div class="widget-title"><h2>Seguridad ciudadana</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="post_list_medium_widget"> 
    <div class="feature-post-list list-post-builder loop-post-content list-with-below-grid ">    
    <div class="image_post feature-item grid_below_image">
                 <a href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/" class="feature-link" title="Alcaldía de Santa Tecla instala 6 cámaras de videovigilancia en bulevar Monseñor Romero">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Alcaldia-Santa-Tecla-e1521673575951-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="post_loop_content">
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:#dd3333" href="http://ultimahora.sv/category/portada/portada-portada/">portada</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67318" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>    
 <h3 class="image-post-title feature_2col"><a href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/">Alcaldía de Santa Tecla instala 6 cámaras de videovigilancia en bulevar Monseñor Romero</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p><p class="post_des">El alcalde de Santa Tecla, Roberto d’Aubuisson, instaló seis nuevas cámaras de videovigilancia en el bulevar Monseñor Arnulfo Romero, esto como parte del proyecto... </p>
<a class="more_button_post" href="http://ultimahora.sv/alcaldia-de-santa-tecla-instala-6-camaras-de-videovigilancia-en-bulevar-monsenor-romero/">Leer más</a>
</div>
 </div>
    </div>



     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow">   
                					
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/concejal-electo-de-chirilagua-fue-asesinado-este-martes/" class="feature-image-link image_post" title="Concejal electo de Chirilagua fue asesinado este martes">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/chirilagua-e1521580818235-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/chirilagua-e1521580818235-100x75.jpg 100w, http://ultimahora.sv/wp-content/uploads/2018/03/chirilagua-e1521580818235-300x224.jpg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/chirilagua-e1521580818235.jpg 484w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/concejal-electo-de-chirilagua-fue-asesinado-este-martes/">Concejal electo de Chirilagua fue asesinado este martes</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/menor-de-edad-es-baleado-por-agente-del-cam-de-santa-tecla/" class="feature-image-link image_post" title="Menor de edad es baleado por agente del CAM de Santa Tecla">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/CAM-NIÑO-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/menor-de-edad-es-baleado-por-agente-del-cam-de-santa-tecla/">Menor de edad es baleado por agente del CAM de Santa Tecla</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/howard-cotto-plantea-hacer-reforma-para-que-medidas-extraordinarias-de-seguridad-sean-permanentes/" class="feature-image-link image_post" title="Howard Cotto plantea hacer reforma para que medidas extraordinarias de seguridad sean permanentes">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Cottito-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/howard-cotto-plantea-hacer-reforma-para-que-medidas-extraordinarias-de-seguridad-sean-permanentes/">Howard Cotto plantea hacer reforma para que medidas extraordinarias de seguridad sean permanentes</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 16, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/pnc-y-fgr-por-cuarta-vez-golpean-finanzas-de-la-ms13/" class="feature-image-link image_post" title="PNC y FGR por cuarta vez golpean finanzas de la MS13">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/detenciones-100x75.jpeg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/detenciones-100x75.jpeg 100w, http://ultimahora.sv/wp-content/uploads/2018/03/detenciones-300x225.jpeg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/detenciones-768x576.jpeg 768w, http://ultimahora.sv/wp-content/uploads/2018/03/detenciones-1024x768.jpeg 1024w, http://ultimahora.sv/wp-content/uploads/2018/03/detenciones.jpeg 1040w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a><a class="post-category-color-text" style="color:" href="http://ultimahora.sv/category/uncategorized/">Uncategorized</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/pnc-y-fgr-por-cuarta-vez-golpean-finanzas-de-la-ms13/">PNC y FGR por cuarta vez golpean finanzas de la MS13</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 16, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/confirman-relanzamiento-de-policia-rural-como-division-de-proteccion-rural/" class="feature-image-link image_post" title="Confirman relanzamiento de Policía Rural como División de Protección Rural">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/1320331-735x400-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#2850ff" href="http://ultimahora.sv/category/arena/">ARENA</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/confirman-relanzamiento-de-policia-rural-como-division-de-proteccion-rural/">Confirman relanzamiento de Policía Rural como División de Protección Rural</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 15, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/la-uca-pide-nuevo-ministro-de-defensa-y-sugiere-que-sea-un-civil/" class="feature-image-link image_post" title="La UCA pide nuevo ministro de Defensa, y sugiere que sea un civil">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/02/tojeira-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2017/02/tojeira-100x75.jpg 100w, http://ultimahora.sv/wp-content/uploads/2017/02/tojeira-300x225.jpg 300w, http://ultimahora.sv/wp-content/uploads/2017/02/tojeira-768x576.jpg 768w, http://ultimahora.sv/wp-content/uploads/2017/02/tojeira.jpg 800w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#8224e3" href="http://ultimahora.sv/category/seguridad-ciudadana/">Seguridad ciudadana</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/la-uca-pide-nuevo-ministro-de-defensa-y-sugiere-que-sea-un-civil/">La UCA pide nuevo ministro de Defensa, y sugiere que sea un civil</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 28, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-5" class="aq-block aq-block-home_large_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-8">
        <div class="widget-title"><h2>Economía</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="post_list_medium_widget"> 
    <div class="feature-post-list list-post-builder loop-post-content list-with-below-grid ">    
    <div class="image_post feature-item grid_below_image">
                 <a href="http://ultimahora.sv/ministro-de-hacienda-impulsara-negociacion-para-consolidar-ley-de-responsabilidad-fiscal/" class="feature-link" title="Ministro de Hacienda impulsará negociación para consolidar Ley de Responsabilidad Fiscal">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Nelson-Fuentes-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="post_loop_content">
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67295" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>    
 <h3 class="image-post-title feature_2col"><a href="http://ultimahora.sv/ministro-de-hacienda-impulsara-negociacion-para-consolidar-ley-de-responsabilidad-fiscal/">Ministro de Hacienda impulsará negociación para consolidar Ley de Responsabilidad Fiscal</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p><p class="post_des">El nuevo ministro de Hacienda, Nelson Fuentes, dijo este miércoles que bajo la actual gestión aún están pendientes las negociaciones para trabajar más en la Ley de... </p>
<a class="more_button_post" href="http://ultimahora.sv/ministro-de-hacienda-impulsara-negociacion-para-consolidar-ley-de-responsabilidad-fiscal/">Leer más</a>
</div>
 </div>
    </div>



     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow">   
                					
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/primer-logro-de-luz-estrella-es-alcanzar-certificacion-para-pupusas-de-olocuilta/" class="feature-image-link image_post" title="Primer logro de Luz Estrella es alcanzar &#8220;certificación&#8221; para pupusas de Olocuilta">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Pupupusas-696x522-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2018/03/Pupupusas-696x522-100x75.jpg 100w, http://ultimahora.sv/wp-content/uploads/2018/03/Pupupusas-696x522-300x225.jpg 300w, http://ultimahora.sv/wp-content/uploads/2018/03/Pupupusas-696x522.jpg 696w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/primer-logro-de-luz-estrella-es-alcanzar-certificacion-para-pupusas-de-olocuilta/">Primer logro de Luz Estrella es alcanzar &#8220;certificación&#8221; para pupusas de Olocuilta</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/monge-no-se-esperan-resultados-sorprendentes-en-economia-con-los-cambios-en-el-gobierno/" class="feature-image-link image_post" title="Monge: No se esperan resultados sorprendentes en economía con los cambios en el Gobierno">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/06/Rigoberto_Monge-e1496411732845-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/monge-no-se-esperan-resultados-sorprendentes-en-economia-con-los-cambios-en-el-gobierno/">Monge: No se esperan resultados sorprendentes en economía con los cambios en el Gobierno</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/el-salvador-recibe-397-8-millones-de-remesas-en-febrero-segun-el-bcr/" class="feature-image-link image_post" title="El Salvador recibe $397.8 millones de remesas en febrero, según el BCR">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/03/Billetes-dolares-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/el-salvador-recibe-397-8-millones-de-remesas-en-febrero-segun-el-bcr/">El Salvador recibe $397.8 millones de remesas en febrero, según el BCR</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 15, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/nuevo-cuscatlan-tendra-modernas-torres-para-complejos-residenciales/" class="feature-image-link image_post" title="Nuevo Cuscatlán tendrá modernas torres para complejos residenciales">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/02/25615548742_34770681a6_b-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/nuevo-cuscatlan-tendra-modernas-torres-para-complejos-residenciales/">Nuevo Cuscatlán tendrá modernas torres para complejos residenciales</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 16, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>									
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/el-salvador-recibio-380-6-millones-en-remesas-en-enero/" class="feature-image-link image_post" title="El Salvador recibió $380.6 millones en remesas en enero">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/04/Dolares-2-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2017/04/Dolares-2-100x75.jpg 100w, http://ultimahora.sv/wp-content/uploads/2017/04/Dolares-2-300x225.jpg 300w, http://ultimahora.sv/wp-content/uploads/2017/04/Dolares-2-768x576.jpg 768w, http://ultimahora.sv/wp-content/uploads/2017/04/Dolares-2.jpg 1024w" sizes="(max-width: 100px) 100vw, 100px" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/el-salvador-recibio-380-6-millones-en-remesas-en-enero/">El Salvador recibió $380.6 millones en remesas en enero</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 14, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 									
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/mas-de-800-turistas-llegaron-este-domingo-a-el-salvador-a-bordo-del-crucero-azamara/" class="feature-image-link image_post" title="Más de 800 turistas llegaron este domingo a El Salvador a bordo del crucero Azamara">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/01/Azamara-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#eeee22" href="http://ultimahora.sv/category/economia/">Economía</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/mas-de-800-turistas-llegaron-este-domingo-a-el-salvador-a-bordo-del-crucero-azamara/">Más de 800 turistas llegaron este domingo a El Salvador a bordo del crucero Azamara</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 28, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-6" class="aq-block aq-block-home_carousel_post aq_span12 aq-first clearfix">        <div class="widget carousel_pagebuilder_wrapper color-4">
        <div class="widget-title"><h2>Negocios</h2></div>		<div class="owl_carousel_builder carousel_pagebuilder">
        
           

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/alcaldia-capitalina-agradece-apertura-de-lecafe-en-el-corazon-del-centro-historico/" class="feature-link" title="Alcaldía capitalina agradece apertura de LeCafe en el corazón del Centro Histórico">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Inauguran-LeCafé-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67188" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/alcaldia-capitalina-agradece-apertura-de-lecafe-en-el-corazon-del-centro-historico/">Alcaldía capitalina agradece apertura de LeCafe en el corazón del Centro Histórico</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 20, 2018</span></p> <p>Los capitalinos podrán deleitar su paladar con una buena taza de café y refrescarse la... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/alcaldia-capitalina-agradece-apertura-de-lecafe-en-el-corazon-del-centro-historico/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                   

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/la-friopack-golden-la-hielea-eco-amigable-para-este-verano/" class="feature-link" title="La “FrioPack Golden” la hielea eco-amigable para este verano">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Screenshot-2018-03-13-at-10.36.53-400x260.png" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="66435" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/la-friopack-golden-la-hielea-eco-amigable-para-este-verano/">La “FrioPack Golden” la hielea eco-amigable para este verano</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 13, 2018</span></p> <p>Golden invita a todos a darle un #refresh a la forma antigua de ver las cosas y le... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/la-friopack-golden-la-hielea-eco-amigable-para-este-verano/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                   

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/proyecto-refresh-la-apuesta-innovadora-de-golden-para-dejar-una-huella-positiva-en-los-salvadorenos/" class="feature-link" title="“Proyecto Refresh“ la apuesta innovadora de Golden para dejar una huella positiva en los salvadoreños">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/02/11-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="64728" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/proyecto-refresh-la-apuesta-innovadora-de-golden-para-dejar-una-huella-positiva-en-los-salvadorenos/">“Proyecto Refresh“ la apuesta innovadora de Golden para dejar una huella positiva en los salvadoreños</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 27, 2018</span></p> <p>Unir a la gente por un mundo mejor, es el sueño de la Constancia, es por es que a... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/proyecto-refresh-la-apuesta-innovadora-de-golden-para-dejar-una-huella-positiva-en-los-salvadorenos/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                   

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/fedecredito-entrega-premios-a-ganadores-de-promocion-gana-facil/" class="feature-link" title="FEDECRÉDITO entrega premios a ganadores de promoción Gana Fácil">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/01/Fedecrédito-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="60907" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/fedecredito-entrega-premios-a-ganadores-de-promocion-gana-facil/">FEDECRÉDITO entrega premios a ganadores de promoción Gana Fácil</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 24, 2018</span></p> <p>Los Bancos de los Trabajadores del Sistema FEDECRÉDITO entregaron a 158 asiduos clientes... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/fedecredito-entrega-premios-a-ganadores-de-promocion-gana-facil/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                   

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/banco-promerica-y-amate-travel-hacen-realidad-tus-vacaciones-sonadas/" class="feature-link" title="Banco Promerica y Amate Travel  hacen realidad tus vacaciones soñadas">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/01/promerica-feria-de-viajes-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="60876" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/banco-promerica-y-amate-travel-hacen-realidad-tus-vacaciones-sonadas/">Banco Promerica y Amate Travel  hacen realidad tus vacaciones soñadas</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 24, 2018</span></p> <p>Banco Promerica y Amate Travel  anunciaron su tradicional feria de viajes... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/banco-promerica-y-amate-travel-hacen-realidad-tus-vacaciones-sonadas/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                   

    <div class="feature-four-column medium-four-columns ">     
    <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/footsolutions-innova-con-atencion-especializada-para-el-cuidado-de-los-pies/" class="feature-link" title="FootSolutions innova con atención especializada para el cuidado de los píes">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2017/12/footsolucion-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#027773" href="http://ultimahora.sv/category/negocios/">Negocios</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="57147" title="Like"><i class="fa fa-heart-o"></i>0</a></div>
</div>
 <h3 class="image-post-title columns_post"><a href="http://ultimahora.sv/footsolutions-innova-con-atencion-especializada-para-el-cuidado-de-los-pies/">FootSolutions innova con atención especializada para el cuidado de los píes</a></h3>      
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Dic 15, 2017</span></p> <p>Electrolab Medic, continúa poniendo a disposición del usuario soluciones integrales... </p>
  <div class="footer_meta"><a href="http://ultimahora.sv/footsolutions-innova-con-atencion-especializada-para-el-cuidado-de-los-pies/" class="footer_meta_readmore">Leer más</a></div>    </div>
         
              
                     
        </div>
        </div>
     
        </div><div id="aq-block-44-7" class="aq-block aq-block-home_large_3main_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-9">
        <div class="widget-title"><h2>Internacionales</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="feature-three-column-home first-child-grid ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/renuncia-presidente-de-peru/" class="feature-link" title="Renuncia presidente de Perú">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/presidente-de-peru-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="67300" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/renuncia-presidente-de-peru/">Renuncia presidente de Perú</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 21, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/renuncia-presidente-de-peru/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
   
	


    <div class="feature-three-column-home ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/quiebra-el-bufete-detras-de-los-panama-papers-mossack-fonseca/" class="feature-link" title="Quiebra el bufete detrás de los Panamá Papers, Mossack Fonseca">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2016/11/1460529024Mossack-Fonseca-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" srcset="http://ultimahora.sv/wp-content/uploads/2016/11/1460529024Mossack-Fonseca-400x260.jpg 400w, http://ultimahora.sv/wp-content/uploads/2016/11/1460529024Mossack-Fonseca-615x400.jpg 615w" sizes="(max-width: 400px) 100vw, 400px" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="66635" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/quiebra-el-bufete-detras-de-los-panama-papers-mossack-fonseca/">Quiebra el bufete detrás de los Panamá Papers, Mossack Fonseca</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 15, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/quiebra-el-bufete-detras-de-los-panama-papers-mossack-fonseca/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
   
	


    <div class="feature-three-column-home ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/smartmatic-ceso-operaciones-en-venezuela/" class="feature-link" title="Smartmatic cesó operaciones en Venezuela">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/000_R64F5-1-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="65740" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/smartmatic-ceso-operaciones-en-venezuela/">Smartmatic cesó operaciones en Venezuela</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 06, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/smartmatic-ceso-operaciones-en-venezuela/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow 3_main_bellow_post_list">   
                 			
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/capturan-a-esposa-del-expresidente-de-honduras-porfirio-lobo/" class="feature-image-link image_post" title="Capturan a esposa del expresidente de Honduras, Porfirio Lobo">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/02/Esposa-Lobo-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/capturan-a-esposa-del-expresidente-de-honduras-porfirio-lobo/">Capturan a esposa del expresidente de Honduras, Porfirio Lobo</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 28, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 				        			
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/oea-pide-a-maduro-no-realizar-elecciones-presidenciales-el-proximo-22-de-abril/" class="feature-image-link image_post" title="OEA pide a Maduro no realizar elecciones presidenciales el próximo 22 de abril">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/02/oea-1-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/oea-pide-a-maduro-no-realizar-elecciones-presidenciales-el-proximo-22-de-abril/">OEA pide a Maduro no realizar elecciones presidenciales el próximo 22 de abril</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 23, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				        			
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/trump-el-salvador-solo-toma-nuestro-dinero/" class="feature-image-link image_post" title="Trump: El Salvador solo toma nuestro dinero">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/08/trump-words-69a90b10-0aa7-11e7-a15f-a58d4a988474-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/trump-el-salvador-solo-toma-nuestro-dinero/">Trump: El Salvador solo toma nuestro dinero</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 23, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 				        			
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/espana-inicia-macrojuicio-en-contra-de-38-miembros-de-la-mara-salvatrucha/" class="feature-image-link image_post" title="España: Inicia “macrojuicio” en contra de 38 miembros de la Mara Salvatrucha">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/02/Salvatrucha-España-770x438-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#dd9933" href="http://ultimahora.sv/category/internacionales/">Internacionales</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/espana-inicia-macrojuicio-en-contra-de-38-miembros-de-la-mara-salvatrucha/">España: Inicia “macrojuicio” en contra de 38 miembros de la Mara Salvatrucha</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-8" class="aq-block aq-block-home_post_right_list_text aq_span12 aq-first clearfix">        <div class="widget main_post_style main_right_post_style_list home_post_right_list_text clearfix color-4">
        <div class="widget-title"><h2>Deportes</h2></div>		<div class="widget_container">
           
<div class="feature-two-column left-post-display-content margin-left-post main-post-right-list  feature-custom">                      
                                <div class="two-content-wrapper main_feature_images main_image_with_list_text">
                    
                <div class="image_post feature-item">
                
                   <a  href="http://ultimahora.sv/fifa-aprueba-uso-del-var-en-rusia-2018/" class="feature-link" title="FIFA aprueba uso del VAR en Rusia 2018">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/var-2-rusia-2018-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
</div>
<div class="main_img_content">
<div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="66828" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/fifa-aprueba-uso-del-var-en-rusia-2018/">FIFA aprueba uso del VAR en Rusia 2018</a></h3>      
 <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 16, 2018</span></p> <p>Fue el mismo presiente de la Federación Internacional de Fútbol Asociado (FIFA), Gianni... </p>
</div>
 
 
    </div>
    </div>
   
 					   <div class="feature-two-column right-post-display-content list-post-right">
                      <ul class="feature-post-list">          
                
                                  
<li class="">
<div class="item-details">
    <span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/barcelona-saca-el-negocio-en-el-campo-del-chelsea/">Barcelona saca el negocio en el campo del Chelsea</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 20, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
            
                               
<li class="">
<div class="item-details">
    <span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/con-pase-filtrado-de-messi-y-gol-de-suarez-inicio-el-gane-del-fc-barcelona/">Con pase filtrado de Messi y gol de Suaréz, inició el gane del FC Barcelona</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 17, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
            
                               
<li class="">
<div class="item-details">
    <span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/el-real-madrid-olvido-lo-que-es-ganar-puntos/">El Real Madrid olvidó lo que es ganar puntos</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Feb 03, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
            
                               
<li class="">
<div class="item-details">
    <span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/alianza-recibe-reconocimiento-de-campeon-en-la-asamblea-legislativa/">Alianza recibe reconocimiento de campeón en la Asamblea Legislativa</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 30, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
            
                               
<li class="">
<div class="item-details">
    <span class="meta-category-small"><a class="post-category-color-text" style="color:#8cffb8" href="http://ultimahora.sv/category/internacionales/deportes/">Deportes</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/fotos-el-magico-recibio-la-elastica-del-cadiz-cf/">FOTOS: El &#8220;Mágico&#8221; recibe la elástica del Cádiz CF</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 29, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
            
                     
			

   </ul>
            </div>
        </div>
         </div>
      
        </div><div id="aq-block-44-9" class="aq-block aq-block-home_large_3main_post_below_list aq_span12 aq-first clearfix">        <div class="widget post_list_medium_widget builder_belowpost color-4">
        <div class="widget-title"><h2>Entretenimiento</h2></div>		<div class="widget_container">
        <div class="post_list_medium">
           
	


    <div class="feature-three-column-home first-child-grid ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/miguel-fortin-deja-a-un-lado-rol-de-analista-para-apoyar-el-talento-de-su-hijo/" class="feature-link" title="Miguel Fortín deja a un lado rol de analista para apoyar el talento de su hijo">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/03/Screenshot-2018-03-16-at-11.54.51-400x260.png" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="66760" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/miguel-fortin-deja-a-un-lado-rol-de-analista-para-apoyar-el-talento-de-su-hijo/">Miguel Fortín deja a un lado rol de analista para apoyar el talento de su hijo</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Mar 16, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/miguel-fortin-deja-a-un-lado-rol-de-analista-para-apoyar-el-talento-de-su-hijo/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
   
	


    <div class="feature-three-column-home ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/generacion-latina-grupo-salsero-salvadoreno-lanza-sencillo-el-son-de-cuscatlan/" class="feature-link" title="Generación Latina, grupo salsero salvadoreño lanza sencillo &#8220;El son de Cuscatlán&#8221;">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/01/generacion-400x260.jpg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="61112" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/generacion-latina-grupo-salsero-salvadoreno-lanza-sencillo-el-son-de-cuscatlan/">Generación Latina, grupo salsero salvadoreño lanza sencillo &#8220;El son de Cuscatlán&#8221;</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 26, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/generacion-latina-grupo-salsero-salvadoreno-lanza-sencillo-el-son-de-cuscatlan/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
   
	


    <div class="feature-three-column-home ">
                    
                <div class="image_post feature-item">
                   <a  href="http://ultimahora.sv/muere-cantante-de-the-craberries/" class="feature-link" title="Muere cantante de The Cranberries">              
<img width="400" height="260" src="http://ultimahora.sv/wp-content/uploads/2018/01/143c01f407ed64a4b3bcbc92d24c05ef80981251-400x260.jpeg" class="attachment-medium-feature size-medium-feature wp-post-image" alt="" /></a>
                     </div>

<div class="wrap_box_style_main feature-custom-below main_post_2col_style">
  <div class="meta_holder">
<span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span><div class="love_this_post_meta"><a href="#" class="jm-post-like" data-post_id="59797" title="Like"><i class="fa fa-heart-o"></i>0</a></div></div>
 <h3 class="image-post-title"><a href="http://ultimahora.sv/muere-cantante-de-the-craberries/">Muere cantante de The Cranberries</a></h3>      
  <p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 15, 2018</span></p>  
 <div class="footer_meta"><a href="http://ultimahora.sv/muere-cantante-de-the-craberries/" class="footer_meta_readmore">Leer más</a></div>   </div>
    </div>

   
     <div class="clear margin-buttons"></div>
      <ul class="feature-post-list large_list_bellow 3_main_bellow_post_list">   
                 			
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/king-flip-si-hubiera-chance-de-entrar-a-la-politica-lo-hago/" class="feature-image-link image_post" title="King Flip: “Si hubiera chance de entrar a la política, lo hago“">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2018/01/Captura-de-pantalla-2018-01-04-a-las-10.16.52-100x75.png" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#1e73be" href="http://ultimahora.sv/category/clase-politica/">Clase política</a><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a><a class="post-category-color-text" style="color:#5b8fbf" href="http://ultimahora.sv/category/lo-ultimo/">Lo último</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/king-flip-si-hubiera-chance-de-entrar-a-la-politica-lo-hago/">King Flip: “Si hubiera chance de entrar a la política, lo hago“</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Ene 04, 2018</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 				        			
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/concurso-canta-con-matices-entrego-1750-dolares-en-premios/" class="feature-image-link image_post" title="Concurso “Canta con Matices“ entregó $1,750 dólares en premios">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/12/DSC03431-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/concurso-canta-con-matices-entrego-1750-dolares-en-premios/">Concurso “Canta con Matices“ entregó $1,750 dólares en premios</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Dic 14, 2017</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				        			
			<li class="large_list_left ">
<a  href="http://ultimahora.sv/steady-rollin-band-lanzara-su-primer-disco-antes-de-fin-de-ano/" class="feature-image-link image_post" title="Steady Rollin Band lanzará su primer disco antes de fin de año">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/12/Rollin-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/steady-rollin-band-lanzara-su-primer-disco-antes-de-fin-de-ano/">Steady Rollin Band lanzará su primer disco antes de fin de año</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Dic 08, 2017</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 				        			
			<li class="large_list_right ">
<a  href="http://ultimahora.sv/fundador-de-espiritu-libre-y-hermano-de-jhosse-lora-muere-atropellado/" class="feature-image-link image_post" title="Fundador de Espíritu Libre y hermano de Jhosse Lora, muere atropellado">              
<img width="100" height="75" src="http://ultimahora.sv/wp-content/uploads/2017/12/fundador-espiritu-libre-100x75.jpg" class="attachment-small-feature size-small-feature wp-post-image" alt="" /></a>
<div class="item-details">
      <span class="meta-category-small"><a class="post-category-color-text" style="color:#c699d8" href="http://ultimahora.sv/category/internacionales/entretenimiento/">Entretenimiento</a></span>
   <h3 class="feature-post-title"><a href="http://ultimahora.sv/fundador-de-espiritu-libre-y-hermano-de-jhosse-lora-muere-atropellado/">Fundador de Espíritu Libre y hermano de Jhosse Lora, muere atropellado</a></h3>
<p class="post-meta meta-main-img"><span class="post-date"><i class="fa fa-clock-o"></i>Dic 05, 2017</span></p>   </div>
   <div class="clearfix"></div>
   </li>
				 <div class="clearfix"></div>				                
         </ul>       
              
                
      </div>
        </div>
        </div>
     
        </div><div id="aq-block-44-10" class="aq-block aq-block-aq_text_block aq_span6 aq-first clearfix"></div></div>
  </div>
  <!-- End content -->
    <!-- Start sidebar -->
<div class="four columns content_display_col3" id="sidebar"><div id="jellywp_fb_likebox_widget-4" class="widget fblikebox_widget">			
<div class="widget_container">   
<div id="fb-root"></div>
<script>(function(d, s, id) {
  var js, fjs = d.getElementsByTagName(s)[0];
  if (d.getElementById(id)) return;
  js = d.createElement(s); js.id = id;
  js.src = "//connect.facebook.net/en_US/all.js#xfbml=1";
  fjs.parentNode.insertBefore(js, fjs);
}(document, 'script', 'facebook-jssdk'));</script>
			

					<div class="fb-like-box" data-href="https://www.facebook.com/ultimahsv/"  data-show-faces="true"  data-stream="true" data-header="true"></div>
	
     <div class="clear"></div>
    </div>
    				

			<div class="margin-bottom"></div></div><div id="text-2" class="widget widget_text">			<div class="textwidget"><a class="twitter-timeline" data-lang="es" data-width="300" data-height="550" data-link-color="#f34035" href="https://twitter.com/ultimahsv"></a> <script async src="//platform.twitter.com/widgets.js" charset="utf-8"></script></div>
		<div class="margin-bottom"></div></div><div id="twitter-follow-2" class="widget widget_twitter-follow"><div class="twitter-follow"><a href="https://twitter.com/intent/follow?screen_name=ultimahsv" class="twitter-follow-button" data-size="large">Seguir a @ultimahsv</a></div><div class="margin-bottom"></div></div></div>  <!-- End sidebar -->
  <div class="clearfix"></div>
  </div>
    
  </div>

<!-- Start footer -->
<footer id="footer-container">

    <div class="footer-columns">
        <div class="row">
                        <div class="four columns"><div id="text-5" class="widget widget_text">			<div class="textwidget"><div style="text-align:center"><img src="http://ultimahora.sv/wp-content/uploads/2016/09/footerlogo.png"></img></div>
<p>Última Hora SV ® 2016</p></div>
		</div></div>
            <div class="four columns"></div>
                                    <div class="four columns"><div id="nav_menu-2" class="widget widget_nav_menu"><div class="menu-footer-container"><ul id="menu-footer" class="menu"><li class="menu-item menu-item-type-post_type menu-item-object-page menu-item-708"><a href="http://ultimahora.sv/contacto/">Contacto</a></li>
</ul></div></div>		<div class="widget">

				
		
			<div class="social_icons_widget">
			<ul class="social-icons-list-widget">
      <li><a href="https://www.facebook.com/ultimahsv" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/facebook.png" alt="Facebook"></a></li>                    <li><a href="https://www.youtube.com/channel/UCxD1dNdPTM7LxkghZ_5wFrA" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/youtube.png" alt="Youtube"></a></li>                         <li><a href="https://twitter.com/ultimahsv" target="_blank"><img src="http://ultimahora.sv/wp-content/themes/nanomag/img/icons/twitter.png" alt="Twitter"></a></li>                                                 </ul> 
			</div>
		</div>
		</div>
     		        </div>
    </div>
          
</footer>
<!-- End footer -->
</div>
<div id="go-top"><a href="#go-top"><i class="fa fa-chevron-up"></i></a></div>
<!-- YouTube Channel 3 --><script type="text/javascript">function ytc_init_MPAU() {jQuery('.ytc-lightbox').magnificPopupAU({disableOn:320,type:'iframe',mainClass:'ytc-mfp-lightbox',removalDelay:160,preloader:false,fixedContentPos:false});}jQuery(window).on('load',function(){ytc_init_MPAU();});jQuery(document).ajaxComplete(function(){ytc_init_MPAU();});</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/f627d.js"></script>

<script type='text/javascript'>
/* <![CDATA[ */
var ajax_var = {"url":"http:\/\/ultimahora.sv\/wp-admin\/admin-ajax.php","nonce":"8cd1c17542"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/4c203.js"></script>

<script type='text/javascript'>
/* <![CDATA[ */
var click_object = {"ajax_url":"http:\/\/ultimahora.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/62f35.js"></script>

<script type='text/javascript'>
/* <![CDATA[ */
var wpcf7 = {"apiSettings":{"root":"http:\/\/ultimahora.sv\/wp-json\/contact-form-7\/v1","namespace":"contact-form-7\/v1"},"recaptcha":{"messages":{"empty":"Por favor, prueba que no eres un robot."}},"cached":"1"};
/* ]]> */
</script>

















<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/9f6c8.js"></script>

<script type='text/javascript'>
/* <![CDATA[ */
var author = {"name":"RU"};
/* ]]> */
</script>
<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/a9198.js"></script>

<script type='text/javascript'>
/* <![CDATA[ */
window.twttr=(function(w){t=w.twttr||{};t._e=[];t.ready=function(f){t._e.push(f);};return t;}(window));
/* ]]> */
</script>
<script type="text/javascript" id="twitter-wjs" async defer src="https://platform.twitter.com/widgets.js" charset="utf-8"></script>

<script type="text/javascript" src="http://ultimahora.sv/wp-content/cache/minify/f394f.js"></script>

</body>
</html>
<!--
Performance optimized by W3 Total Cache. Learn more: https://www.w3-edge.com/products/

Almacenamiento en caché de objetos 7840/117 objetos que utilizan disk
Page Caching using disk: enhanced (Page is front page) 
Red de Entrega de Contenido vía N/A
Minificado usando disk
Caching de base de datos 28/219 consultas en 0.150 segundos usando disk

Served from: ultimahora.sv @ 2018-03-22 04:05:33 by W3 Total Cache
-->