
<!DOCTYPE html>
<html xmlns="http://www.w3.org/1999/xhtml" xml:lang="es-es" lang="es-es" dir="ltr">
<head>

    <meta name="viewport" content="width=device-width, initial-scale=1.0">

  <base href="http://fdim.org.sv/" />
  <meta http-equiv="content-type" content="text/html; charset=utf-8" />
  <meta name="keywords" content="FDIM, federación democrática internacional de mujeres, federación mundial de mujeres" />
  <meta name="description" content="Federación Democrática Internacional de Mujeres" />
  <meta name="generator" content="Joomla! - Open Source Content Management" />
  <title>FDIM - FDIM | Federación Democrática Internacional de Mujeres</title>
  <link href="http://fdim.org.sv/?view=featured" rel="canonical" />
  <link href="/index.php?format=feed&amp;type=rss" rel="alternate" type="application/rss+xml" title="RSS 2.0" />
  <link href="/index.php?format=feed&amp;type=atom" rel="alternate" type="application/atom+xml" title="Atom 1.0" />
  <link href="/templates/it_community2/favicon.ico" rel="shortcut icon" type="image/vnd.microsoft.icon" />
  <link href="http://fdim.org.sv/index.php/component/search/?format=opensearch" rel="search" title="Buscar FDIM" type="application/opensearchdescription+xml" />
  <link rel="stylesheet" href="/plugins/system/iceshortcodes/assets/iceshortcodes.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/bootstrap/css/bootstrap.min.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/font-awesome/css/font-awesome.min.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/bootstrap/css/bootstrap-responsive.min.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/css/joomla.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/css/modules.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/css/general.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/css/pages.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/css/responsive.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_djimageslider/themes/default/css/djimageslider.css" type="text/css" />
  <link rel="stylesheet" href="/media/djextensions/magnific/magnific.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_featured_youtube_slider/css/style-responsive.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_fblikeboxslider/css/style.css" type="text/css" />
  <link rel="stylesheet" href="/modules/mod_iceslideshow/assets/style.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/html/mod_icemegamenu/css/default_icemegamenu.css" type="text/css" />
  <link rel="stylesheet" href="/templates/it_community2/html/mod_icemegamenu/css/default_icemegamenu-reponsive.css" type="text/css" />
  <style type="text/css">

	.responsive.modfytslider{
		background: #d9d9d9;
	}
	
	.responsive .sliderwrapper{
		background: #d9d9d9;
	}
	
	.responsive .sliderwrapper .contentdiv{
		background: #ffffff;
	}

	.responsive .paginationfytslide{
		background: #cccccc;
	}
	
	.responsive .paginationfytslide a img,.paginationfytslide a:visited img{
		background: #d9d9d9;
	}
	
	.responsive .paginationfytslide a:hover img{
		background: #cccccc;
	}
	
	@media screen and (min-width: 378px) and (max-width: 470px){
		.responsive .paginationfytslide-inner a img,
		.responsive .paginationfytslide-inner img{
			width:22%!important;
		}
	}
	
	@media screen and (min-width: 471px) and (max-width: 780px){
		.responsive .paginationfytslide-inner a img,
		.responsive .paginationfytslide-inner img{
			width:22%!important;
		}
	}
	
	@media screen and (min-width: 781px) and (max-width: 991px){
		.responsive .paginationfytslide-inner a img,
		.responsive .paginationfytslide-inner img{
			width:47%!important;
		}
	}

#goog-gt-tt {display:none !important;}
.goog-te-banner-frame {display:none !important;}
.goog-te-menu-value:hover {text-decoration:none !important;}
body {top:0 !important;}
#google_translate_element2 {display:none!important;}

        a.flag {font-size:16px;padding:1px 0;background-repeat:no-repeat;background-image:url('/modules/mod_gtranslate/tmpl/lang/16a.png');}
        a.flag:hover {background-image:url('/modules/mod_gtranslate/tmpl/lang/16.png');}
        a.flag img {border:0;}
        a.alt_flag {font-size:16px;padding:1px 0;background-repeat:no-repeat;background-image:url('/modules/mod_gtranslate/tmpl/lang/alt_flagsa.png');}
        a.alt_flag:hover {background-image:url('/modules/mod_gtranslate/tmpl/lang/alt_flags.png');}
        a.alt_flag img {border:0;}
    
  </style>
  <script src="/media/system/js/mootools-core.js" type="text/javascript"></script>
  <script src="/media/system/js/core.js" type="text/javascript"></script>
  <script src="/media/system/js/caption.js" type="text/javascript"></script>
  <script src="/media/jui/js/jquery.min.js" type="text/javascript"></script>
  <script src="/media/jui/js/jquery-noconflict.js" type="text/javascript"></script>
  <script src="/templates/it_community2/bootstrap/js/bootstrap.min.js" type="text/javascript"></script>
  <script src="/media/djextensions/jquery-easing/jquery.easing.min.js" type="text/javascript" defer="defer"></script>
  <script src="/modules/mod_djimageslider/assets/js/slider.js?v=" type="text/javascript" defer="defer"></script>
  <script src="/media/djextensions/magnific/magnific.js" type="text/javascript" defer="defer"></script>
  <script src="/modules/mod_djimageslider/assets/js/magnific-init.js" type="text/javascript" defer="defer"></script>
  <script src="/modules/mod_featured_youtube_slider/library/contentslider.js" type="text/javascript"></script>
  <script type="text/javascript">
window.addEvent('load', function() {
				new JCaption('img.caption');
			});
    jQuery(document).ready(function(){ 
			
			 jQuery(window).scroll(function(){
				if ( jQuery(this).scrollTop() > 1000) {
					 jQuery('#gotop').addClass('gotop_active');
				} else {
					 jQuery('#gotop').removeClass('gotop_active');
				}
			}); 
			
			jQuery('.scrollup').click(function(){
				jQuery("html, body").animate({ scrollTop: 0 }, 600);
				return false;
			});
			
 
		});

jQuery(document).ready(function(){ 
		
	if (jQuery('body').height() > 1200) {
		 jQuery('body').addClass('body_effect_bottom');
	}
	
	jQuery( "#cGallery .photoLoad" ).append( '<ul class="ice_css3_loading"><li></li><li></li><li></li><li></li></ul>' );
	
	jQuery("[rel='tooltip']").tooltip();
	
	
	jQuery("#language img").hover(function () {
		jQuery("#language img").css({opacity : .25});
	  }, 
	  function () {
		jQuery("#language img").css({ opacity : 1});
	  }
	);	
	
});

	jQuery(document).ready(function() {     
	jQuery('.mainmenu').hover(function(){     
		jQuery('#iceslideshow > div > div:first-child').addClass('icemegamenu-hover');    
	},     
	function(){    
	   jQuery('#iceslideshow > div > div:first-child').removeClass('icemegamenu-hover');     
	});
	});   

if (("ontouchstart" in document.documentElement)) {
	document.documentElement.className += "with-touch";
}else {
	document.documentElement.className += "no-touch";
}
				

  </script>
  <script type="text/javascript" src="http://s7.addthis.com/js/300/addthis_widget.js"></script>


	<style type="text/css" media="screen">

	
/* Sidebar is "left" */
#middlecol { float:right !important;}


/* Custom CSS code throught paramters */
</style>

<!-- Template Styles  -->
<link id="stylesheet" rel="stylesheet" type="text/css" href="/templates/it_community2/css/styles/style1.css" />

<!-- Resposnive Template Styles -->
<link id="stylesheet-responsive" rel="stylesheet" type="text/css" href="/templates/it_community2/css/styles/style1_responsive.css" />



<!-- Google Fonts -->
<link href='http://fonts.googleapis.com/css?family=Rosario|Open+Sans|Coming+Soon' rel='stylesheet' type='text/css' />

<!--[if lte IE 8]>
<link rel="stylesheet" type="text/css" href="/templates/it_community2/css/ie8.css" />
<script src="/templates/it_community2/js/respond.min.js"></script>
<![endif]-->

<!--[if lt IE 9]>
    <script src="/media/jui/js/html5.js"></script>
<![endif]-->


<!--[if !IE]><!-->
<script>  
if(Function('/*@cc_on return document.documentMode===10@*/')()){
    document.documentElement.className+=' ie10';
}
</script>
<!--<![endif]-->  

<style type="text/css">

/* IE10 hacks. add .ie10 before */
.ie10 ul#ice-switcher {
	padding-right:20px;}  
	.ie10 ul#ice-switcher:hover {
		padding-right:35px}

.ie10 ul#ice-switcher li.active a,
.ie10 ul#ice-switcher li a:hover {
	padding-top:0;
	padding-bottom:0}
					
.ie10 ul#ice-switcher li a span {
	padding-left:30px;}
	
.ie10 #gotop .scrollup {
	right:40px;}

</style>




        
</head>

<body class="">   

    <!-- header -->
    <header id="header" class="container">
    
        <div id="logo">	
        	<a href="/"><img class="logo" src="http://fdim.org.sv/images/sampledata/icetheme/logo.png" alt="FDIM" /></a>	
        </div>
            
                <div id="language">	
           

<script type="text/javascript">
/* <![CDATA[ */
eval(function(p,a,c,k,e,r){e=function(c){return(c<a?'':e(parseInt(c/a)))+((c=c%a)>35?String.fromCharCode(c+29):c.toString(36))};if(!''.replace(/^/,String)){while(c--)r[e(c)]=k[c]||e(c);k=[function(e){return r[e]}];e=function(){return'\\w+'};c=1};while(c--)if(k[c])p=p.replace(new RegExp('\\b'+e(c)+'\\b','g'),k[c]);return p}('6 7(a,b){n{4(2.9){3 c=2.9("o");c.p(b,f,f);a.q(c)}g{3 c=2.r();a.s(\'t\'+b,c)}}u(e){}}6 h(a){4(a.8)a=a.8;4(a==\'\')v;3 b=a.w(\'|\')[1];3 c;3 d=2.x(\'y\');z(3 i=0;i<d.5;i++)4(d[i].A==\'B-C-D\')c=d[i];4(2.j(\'k\')==E||2.j(\'k\').l.5==0||c.5==0||c.l.5==0){F(6(){h(a)},G)}g{c.8=b;7(c,\'m\');7(c,\'m\')}}',43,43,'||document|var|if|length|function|GTranslateFireEvent|value|createEvent||||||true|else|doGTranslate||getElementById|google_translate_element2|innerHTML|change|try|HTMLEvents|initEvent|dispatchEvent|createEventObject|fireEvent|on|catch|return|split|getElementsByTagName|select|for|className|goog|te|combo|null|setTimeout|500'.split('|'),0,{}))
/* ]]> */
</script>


<div id="google_translate_element2"></div>
<script type="text/javascript">function googleTranslateElementInit2() {new google.translate.TranslateElement({pageLanguage: 'es', autoDisplay: false}, 'google_translate_element2');}</script>
<script type="text/javascript" src="//translate.google.com/translate_a/element.js?cb=googleTranslateElementInit2"></script>

<a href="#" onclick="doGTranslate('es|es');return false;" title="Spanish" class="flag nturl" style="background-position:-600px -200px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="16" width="16" alt="Spanish" /></a> <a href="#" onclick="doGTranslate('es|en');return false;" title="English" class="alt_flag" style="background-position:-0px -0px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="16" width="16" alt="English" /></a>  <a href="#" onclick="doGTranslate('es|fr');return false;" title="French" class="flag nturl" style="background-position:-200px -100px;"><img src="/modules/mod_gtranslate/tmpl/lang/blank.png" height="16" width="16" alt="French" /></a> 
        </div> 
                
                <div id="search">
            <div class="search">
    <form action="/index.php" method="post" class="form-inline">
    		<label for="mod-search-searchword" class="element-invisible">Buscar...</label> <input name="searchword" id="mod-search-searchword" maxlength="20"  class="inputbox search-query" type="text" size="20" value="Buscar..."  onblur="if (this.value=='') this.value='Buscar...';" onfocus="if (this.value=='Buscar...') this.value='';" /> <button class="button btn btn-primary" onclick="this.form.searchword.focus();">Go</button>    	<input type="hidden" name="task" value="search" />
    	<input type="hidden" name="option" value="com_search" />
    	<input type="hidden" name="Itemid" value="435" />
    </form>
</div>

        </div>
          
        
                
        <div id="mainmenu" class="clearfix">
            <div class="mainmenu">
                <div class="icemegamenu"><div class="ice-megamenu-toggle"><a data-toggle="collapse" data-target=".nav-collapse" href="#">Menu</a></div><div class="nav-collapse icemegamenu collapse"><ul id="icemegamenu" class="meganizr mzr-slide mzr-responsive"><li id="iceMenu_435" class="iceMenuLiLevel_1 active"><a href="http://fdim.org.sv/" class="icemega_active iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Inicio</span></a></li><li id="iceMenu_475" class="iceMenuLiLevel_1 mzr-drop parent"><a class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Presidencia</span></a><ul class="icesubMenu icemodules sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_476" class="iceMenuLiLevel_2"><a href="/index.php/presidencia/biografia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Biografía</span></a></li><li id="iceMenu_749" class="iceMenuLiLevel_2"><a href="/index.php/presidencia/vice-presidencia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Secretariado Mundial</span></a></li></ul></div></li></ul></li><li id="iceMenu_750" class="iceMenuLiLevel_1 mzr-drop parent"><a class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Conócenos</span></a><ul class="icesubMenu icemodules sub_level_1" style="width:280px"><li><div style="float:left;width:280px" class="iceCols"><ul><li id="iceMenu_477" class="iceMenuLiLevel_2"><a href="/index.php/conocenos/historia" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Historia</span></a></li><li id="iceMenu_810" class="iceMenuLiLevel_2"><a href="/index.php/conocenos/estructura" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Estructura</span></a></li><li id="iceMenu_811" class="iceMenuLiLevel_2"><a href="/index.php/conocenos/xvi-congreso-fdim" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">XVI Congreso FDIM</span></a></li></ul></div></li></ul></li><li id="iceMenu_540" class="iceMenuLiLevel_1 mzr-drop parent"><a class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Regiones</span></a><ul class="icesubMenu icemodules sub_level_1" style="width:300px"><li><div style="float:left;width:300px" class="iceCols"><ul><li id="iceMenu_745" class="iceMenuLiLevel_2"><a href="/index.php?Itemid=745" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Asia</span></a></li><li id="iceMenu_746" class="iceMenuLiLevel_2"><a href="/index.php/regiones/america-y-el-caribe" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">América y El Caribe</span></a></li><li id="iceMenu_747" class="iceMenuLiLevel_2"><a href="/index.php/regiones/europa" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Europa</span></a></li><li id="iceMenu_748" class="iceMenuLiLevel_2"><a href="/index.php/regiones/africa" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">África</span></a></li><li id="iceMenu_791" class="iceMenuLiLevel_2"><a href="/index.php/regiones/paises-arabes" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Países Árabes</span></a></li></ul></div></li></ul></li><li id="iceMenu_807" class="iceMenuLiLevel_1"><a href="/index.php/noticias" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Noticias</span></a></li><li id="iceMenu_808" class="iceMenuLiLevel_1"><a href="/index.php/comunicados" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Comunicados</span></a></li><li id="iceMenu_809" class="iceMenuLiLevel_1"><a href="/index.php/publicaciones" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Publicaciones</span></a></li><li id="iceMenu_798" class="iceMenuLiLevel_1"><a href="http://fdim.org.sv/webmail" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Correo</span></a></li><li id="iceMenu_661" class="iceMenuLiLevel_1"><a href="/index.php/contactenos" class=" iceMenuTitle"><span class="icemega_title icemega_nosubtitle">Contáctenos</span></a></li></ul></div></div>
<script type="text/javascript">
	jQuery(document).ready(function(){
		var browser_width1 = jQuery(window).width();
		jQuery("#icemegamenu").find(".icesubMenu").each(function(index){
			var offset1 = jQuery(this).offset();
			var xwidth1 = offset1.left + jQuery(this).width();
			if(xwidth1 >= browser_width1){
				jQuery(this).addClass("ice_righttoleft");
			}
		});
		
	})
	jQuery(window).resize(function() {
		var browser_width = jQuery(window).width();
		jQuery("#icemegamenu").find(".icesubMenu").removeClass("ice_righttoleft");
		jQuery("#icemegamenu").find(".icesubMenu").each(function(index){
			var offset = jQuery(this).offset();
			var xwidth = offset.left + jQuery(this).width();
			
			if(xwidth >= browser_width){
				jQuery(this).addClass("ice_righttoleft");
			}
		});
	});
</script>
            </div>
        </div>

		        <div id="iceslideshow">
            
<div id="iceslideshow366" class="iceslideshow carousel slide Slide Next carousel-fade mootools-noconflict">
       
	<div id="ice_slideshow_preload366" class="ice_preload">
    	
         <div id="movingBallG">
			<div class="movingBallLineG">
			</div>
            <div id="movingBallG_1" class="movingBallG">
            </div>
		</div>
    
    </div>
        
        <div class="carousel-inner">
								<div class="item active">
					
					<img src="http://fdim.org.sv/images/icethumbs/1170x420/100/images/image24.jpg" title="item4" alt="item4" width="1170px" height="420px" />	
						
							
						
							<div class="carousel-caption">
                              
							                              <div class="mod-description">
                              	
                                 
                                  
                              </div>
                                                        
														  
							</div>
							
												
					  </div>
										<div class="item ">
					
					<img src="http://fdim.org.sv/images/icethumbs/1170x420/100/images/image02.jpg" title="item2" alt="item2" width="1170px" height="420px" />	
						
							
						
							<div class="carousel-caption">
                              
							                              <div class="mod-description">
                              	
                                 
                                  
                              </div>
                                                        
														  
							</div>
							
												
					  </div>
										<div class="item ">
					
					<img src="http://fdim.org.sv/images/icethumbs/1170x420/100/images/image03.jpg" title="item3" alt="item3" width="1170px" height="420px" />	
						
							
						
							<div class="carousel-caption">
                              
							                              <div class="mod-description">
                              	
                                 
                                  
                              </div>
                                                        
														  
							</div>
							
												
					  </div>
					        </div><!-- .carousel-inner -->
					<!--  next and previous controls here
				  href values must reference the id for this carousel -->
             <div class="iceslideshow_arrow">
			  <a class="carousel-control left" href="#iceslideshow366" data-slide="prev">&lsaquo;</a>
			  <a class="carousel-control right" href="#iceslideshow366" data-slide="next">&rsaquo;</a>
              </div>
		</div>

<script type="text/javascript">
	jQuery(window).load (function () { 
	  jQuery('#ice_slideshow_preload366').removeClass('ice_preload')
	});
</script>



    
<script type="text/javascript">

if (typeof jQuery != 'undefined') { 
	(function($) { 
		$(document).ready(function(){
			$('.carousel').each(function(index, element) {
			$(this)[index].slide = null;
			});
		});
	})(jQuery);
}

jQuery(document).ready(function(){

	jQuery('#iceslideshow366').carousel(
	
		{ interval: 5000, pause:"hover" }
		
	
	);
});
	  
</script>


        </div>
                
	</header><!-- /header -->


	    <div id="services" class="container">
        

<div class="custom"  >
	<div class="row">
<div class="span3"><img src="/images/SERVICES/Maria_Lisa_Cinciari_Rodano.jpg" alt="Maria Lisa Cinciari Rodano" width="129" height="64" />
<h3>Maria Lisa Cinciari</h3>
<p>"Con la fundaci&oacute;n de la FDIM teniamos la esperanza de aportar a construir un nuevo mundo y la conquista plena de los derechos de las mujeres"</p>
</div>
<div class="span3"><img src="/images/SERVICES/Linda_Matar.png" alt="Linda Matar" width="129" height="115" />
<h3>Linda Matar</h3>
<p>"Seguiremos demostrando que los sue&ntilde;os no se miden por la edad, estos contin&uacute;an mientras haya un coraz&oacute;n latiendo"</p>
</div>
<div class="span3"><img src="/images/photo4.jpg" alt="Sample Photo" width="150" height="150" />
<h3>Melida Anaya Montes</h3>
<p>"En los momentos mas dificiles hay que tener la mente fria y el corazon ardiente de amor por la poblacion"</p>
</div>
<div class="span3"><img src="/images/photo6.jpg" alt="Sample Photo" width="150" height="150" />
<h3>Vilma Esp&iacute;n</h3>
<p>"Una gran maestra de la vida, distinguida por su amor y de dedicaci&oacute;n a la obra de la revoluci&oacute;n"</p>
</div>
</div></div>

    </div>
    

	<!-- content -->
	<section id="content" class="container">

		<div class="newsflash">
</div>



 <script src="http://code.jquery.com/jquery-latest.js"></script>

	<style type="text/css">
#on {
  visibility: visible;
}
#off {
  visibility: hidden;
}
#facebook_div {
  width: 196px;
  height: 340px;
  overflow: hidden;
}
#twitter_div {
  width: 276px;
  height: 280px;
  overflow: hidden;
}
#NBT_div {
  width: 300px;
  height: 97px;
  overflow: hidden;
}
/* right side style */
#twitter_right {
  z-index: 10004;
  border: 2px solid #6CC5FF;
  background-color: #6CC5FF;
  width: 246px;
  height: 280px;
  position: fixed;
  right: -250px;
}
#twitter_right_img {
  position: absolute;
  top: -2px;
  left: -35px;
  border: 0;
}
#NBT_right {
  z-index: 10003;
  border: 2px solid #303030;
  background-color: #fff;
  width: 300px;
  height: 97px;
  position: fixed;
}
#NBT_right img {
  position: absolute;
  top: -2px;
  left: -101px;
}
/* left side style */
#twitter_left {
  z-index: 10004;
  border: 2px solid #6CC5FF;
  background-color: #6CC5FF;
  width: 246px;
  height: 280px;
  position: fixed;
  left: -250px;
}
#twitter_left_img {
  position: absolute;
  top: -2px;
  right: -35px;
  border: 0;
}

</style>
<script type="text/javascript">

jQuery(document).ready(function () {
  jQuery("#twitter_right").hover(function () {
    jQuery(this).stop(true, false).animate({
      right: 0
    }, 500);
  }, function () {
    jQuery("#twitter_right").stop(true, false).animate({
      right: -250
    }, 500);
  });
  
});
</script>
<div id="twitter_right" style="top: 250px;">
 <div id="twitter_div">
		<img id="twitter_right_img" src="http://fdim.org.sv/modules/mod_twitterslider/twitter_right.png" />
 	
		<div id="twitterfanbox">
<a class="twitter-timeline" data-link-color="#f5784f" data-theme="light" data-chrome=""   href="https://twitter.com/@fdim_" width="246" height="280">Tweets by @@fdim_</a>

<script async src="//platform.twitter.com/widgets.js" charset="utf-8"></script>		</div>
		
	</div>
	<div style="font-size: 9px; color: #808080; font-weight: normal; font-family: tahoma,verdana,arial,sans-serif; line-height: 1.28; text-align: right; direction: ltr;"><a class="nolink"></a></div>
</div>
	

	<div id="awesome_facebook">
        <div id="facebookbox1"
        
                    <div style="right: -310px; top: 110px; z-index: 10000;">
                    <div id="facebookbox2" style="text-align: left;height:px;">
            
                  
                <img style="top: 0px;left:-46px;" src="/modules/mod_fblikeboxslider/images/fb.png" alt="">
                
               
            <div id="fb-root"></div>
      <script>
        (function(d, s, id) {
          var js, fjs = d.getElementsByTagName(s)[0];
          if (d.getElementById(id)) return;
          js = d.createElement(s); js.id = id;
          js.src = "//connect.facebook.net/en_US/sdk.js#xfbml=1&version=v2.0";
          fjs.parentNode.insertBefore(js, fjs);
        }(document, 'script', 'facebook-jssdk'));
            </script>  
            <div class="fb-like-box" data-href="https://www.facebook.com/federaciondemocraticainternacionaldemujeres" data-colorscheme="light"  
              data-show-faces="true"   data-header="yes"  
             data-width="300"  data-height="350"
               data-stream="true"                data-show-border="true">             </div>
            
            <div style="font-size: 9px; color: #808080; font-weight: normal; font-family: tahoma,verdana,arial,sans-serif; line-height: 1.28; text-align: right; direction: ltr;"><a class="nolink"></a></div>

            
         </div>


        </div>
        
    </div>
  
  <script type="text/javascript">
    jQuery.noConflict();
    jQuery(function (){
    jQuery(document).ready(function()
    {
    jQuery.noConflict();
    jQuery(function (){
    jQuery("#facebookbox1").hover(function(){ 
    jQuery('#facebookbox1').css('z-index',101009);
    
        
    jQuery(this).stop(true,false).animate({right:  0}, 500); },
    function(){ 
    jQuery('#facebookbox1').css('z-index',10000);
    jQuery("#facebookbox1").stop(true,false).animate({right: -310}, 500); });
    });}); });
    
    </script>


    
    	         
         
        <!-- promo --> 
		        
          
		<div class="row">
        
            <!-- Middle Col -->
            <div id="middlecol" class="span8">
            
                <div class="inside">
                                           
                    
<div id="system-message-container">
<div id="system-message">
</div>
</div>
                
                    <div class="blog-featured">

	
		
		<div class="items-row cols-1 row-0 row-fluid">
					<div class="item column-1 span12">
			

	<h2 class="item-title">
			<a href="/index.php/38-uncategorised/noticias/210-lucha-asesinato-y-racismo-estructural"> Lucha, asesinato y racismo estructural</a>
		</h2>




	<dl class="article-info  muted">
		<dt class="article-info-term">
		Detalles		</dt>

		
		
		
		
					
			
							<dd class="hits">
					<span class="icon-eye-open"></span>
					Visto: 117				</dd>
			
			</dl>

		<div class="pull-left item-image"> <img
		src="/images/MARIELLE.png" alt=""/> </div>

	 <p>&nbsp;</p>
<p style="text-align: center;"><em><em style="text-align: center;">Tras el asesinato de Marielle Franco, el Foro Social Mundial se moviliz&oacute; para exigir justicia por el crimen de la militante feminista y de derechos humanos. La responsabilidad del Gobierno, la violencia contra las mujeres, racismo y el genocidio negro.</em></em></p>
 <div class='joomla_add_this'><!-- AddThis Button BEGIN -->
<script type='text/javascript'>
var addthis_product = 'jlp-2.0';
var addthis_config = {
pubid:'ra-51cd8ef9387066c4',
ui_hover_direction:false,
data_track_clickback:true,
ui_language:'en',
ui_use_css:true
}
</script>
<div class="addthis_toolbox addthis_default_style " addthis:url='http://fdim.org.sv/index.php/38-uncategorised/noticias/210-lucha-asesinato-y-racismo-estructural' addthis:title='Lucha, asesinato y racismo estructural'>
									<a class="addthis_button_preferred_1"></a>
									<a class="addthis_button_preferred_2"></a>
									<a class="addthis_button_preferred_3"></a>
									<a class="addthis_button_preferred_4"></a>
									<a class="addthis_button_compact"></a>
									<a class="addthis_counter addthis_bubble_style"></a>
								</div><!-- AddThis Button END -->
</div>


	<p class="readmore"><a class="btn" href="/index.php/38-uncategorised/noticias/210-lucha-asesinato-y-racismo-estructural"> <span class="icon-chevron-right"></span>

	Leer más...
	</a></p>



			</div>
			
			
		</div>
		
	
		
		<div class="items-row cols-1 row-1 row-fluid">
					<div class="item column-1 span12">
			

	<h2 class="item-title">
			<a href="/index.php/38-uncategorised/noticias/209-farc-resultados-electorales-reafirman-necesidad-de-avanzar-hacia-una-reforma-politico-electoral-de-caracter-estructural"> FARC: Resultados electorales reafirman necesidad de avanzar hacia una reforma político-electoral de carácter estructural.</a>
		</h2>




	<dl class="article-info  muted">
		<dt class="article-info-term">
		Detalles		</dt>

		
		
		
		
					
			
							<dd class="hits">
					<span class="icon-eye-open"></span>
					Visto: 65				</dd>
			
			</dl>

		<div class="pull-left item-image"> <img
		src="/images/colombia.png" alt=""/> </div>

	 <p><span style="text-align: center;"><span style="text-align: justify;">Fuerza Alternativa Revolucionaria del Com&uacute;n (FARC) declar&oacute; en un comunicado de prensa que los resultados electorales del 11 de marzo no modificaron de manera esencial la estructura del Congreso de la Rep&uacute;blica.&nbsp;</span></span></p>
 <div class='joomla_add_this'><!-- AddThis Button BEGIN -->
<script type='text/javascript'>
var addthis_product = 'jlp-2.0';
var addthis_config = {
pubid:'ra-51cd8ef9387066c4',
ui_hover_direction:false,
data_track_clickback:true,
ui_language:'en',
ui_use_css:true
}
</script>
<div class="addthis_toolbox addthis_default_style " addthis:url='http://fdim.org.sv/index.php/38-uncategorised/noticias/209-farc-resultados-electorales-reafirman-necesidad-de-avanzar-hacia-una-reforma-politico-electoral-de-caracter-estructural' addthis:title='FARC: Resultados electorales reafirman necesidad de avanzar hacia una reforma político-electoral de carácter estructural.'>
									<a class="addthis_button_preferred_1"></a>
									<a class="addthis_button_preferred_2"></a>
									<a class="addthis_button_preferred_3"></a>
									<a class="addthis_button_preferred_4"></a>
									<a class="addthis_button_compact"></a>
									<a class="addthis_counter addthis_bubble_style"></a>
								</div><!-- AddThis Button END -->
</div>


	<p class="readmore"><a class="btn" href="/index.php/38-uncategorised/noticias/209-farc-resultados-electorales-reafirman-necesidad-de-avanzar-hacia-una-reforma-politico-electoral-de-caracter-estructural"> <span class="icon-chevron-right"></span>

	Leer más...
	</a></p>



			</div>
			
			
		</div>
		
	
		
		<div class="items-row cols-1 row-2 row-fluid">
					<div class="item column-1 span12">
			

	<h2 class="item-title">
			<a href="/index.php/38-uncategorised/noticias/208-llaman-a-instalar-tribunal-de-los-pueblos-sobre-los-crimenes-de-estados-unidos-contra-puerto-rico"> Llaman a instalar Tribunal de los pueblos sobre los crímenes de Estados Unidos contra Puerto Rico</a>
		</h2>




	<dl class="article-info  muted">
		<dt class="article-info-term">
		Detalles		</dt>

		
		
		
		
					
			
							<dd class="hits">
					<span class="icon-eye-open"></span>
					Visto: 307				</dd>
			
			</dl>

		<div class="pull-left item-image"> <img
		src="/images/puerto-rico libre.png" alt=""/> </div>

	 <p>El Tribunal se estar&iacute;a instalando el &uacute;ltimo s&aacute;bado de octubre de 2018 para exponer la responsabilidad de EUA en el cometido de m&uacute;ltiples violaciones contra el pueblo boricua durante los 120 a&ntilde;os de invasi&oacute;n y ocupaci&oacute;n.</p>
 <div class='joomla_add_this'><!-- AddThis Button BEGIN -->
<script type='text/javascript'>
var addthis_product = 'jlp-2.0';
var addthis_config = {
pubid:'ra-51cd8ef9387066c4',
ui_hover_direction:false,
data_track_clickback:true,
ui_language:'en',
ui_use_css:true
}
</script>
<div class="addthis_toolbox addthis_default_style " addthis:url='http://fdim.org.sv/index.php/38-uncategorised/noticias/208-llaman-a-instalar-tribunal-de-los-pueblos-sobre-los-crimenes-de-estados-unidos-contra-puerto-rico' addthis:title='Llaman a instalar Tribunal de los pueblos sobre los crímenes de Estados Unidos contra Puerto Rico'>
									<a class="addthis_button_preferred_1"></a>
									<a class="addthis_button_preferred_2"></a>
									<a class="addthis_button_preferred_3"></a>
									<a class="addthis_button_preferred_4"></a>
									<a class="addthis_button_compact"></a>
									<a class="addthis_counter addthis_bubble_style"></a>
								</div><!-- AddThis Button END -->
</div>


	<p class="readmore"><a class="btn" href="/index.php/38-uncategorised/noticias/208-llaman-a-instalar-tribunal-de-los-pueblos-sobre-los-crimenes-de-estados-unidos-contra-puerto-rico"> <span class="icon-chevron-right"></span>

	Leer más...
	</a></p>



			</div>
			
			
		</div>
		
	

	<div class="pagination">

					<p class="counter pull-right">
				Página 1 de 29			</p>
						<ul class="pagination-list"><li class="disabled"><a><i class="icon-first"></i></a></li><li class="disabled"><a><i class="icon-previous"></i></a></li><li class="active"><a>1</a></li><li><a title="2" href="/index.php?start=3" class="pagenav">2</a><li><li><a title="3" href="/index.php?start=6" class="pagenav">3</a><li><li><a title="4" href="/index.php?start=9" class="pagenav">4</a><li><li><a title="5" href="/index.php?start=12" class="pagenav">...</a><li><li><a title="6" href="/index.php?start=15" class="pagenav">6</a><li><li><a title="7" href="/index.php?start=18" class="pagenav">7</a><li><li><a title="8" href="/index.php?start=21" class="pagenav">8</a><li><li><a title="9" href="/index.php?start=24" class="pagenav">9</a><li><li><a title="10" href="/index.php?start=27" class="pagenav">10</a><li><li><a title="Siguiente" href="/index.php?start=3" class="pagenav">Siguiente</a><li><li><a title="Final" href="/index.php?start=84" class="pagenav">Final</a><li></ul>	</div>

</div>

                
                </div>
            
            </div>
            <!-- / Middle Col  -->
                
			  
            <!-- sidebar -->
            <div id="sidebar" class="span4 " >
                <div class="inside">    
                    		
		<div class="sidebar_module sidebar_module_">
        	
			                    <h3 class="sidebar_module_heading"><span>Zona Multimedia</span></h3>
                			
           
                <div class="sidebar_module_content"><div class="responsive modfytslider">
<div id="fytslider380" class="sliderwrapper">
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/dYqQQ8k8ETs?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/rGrPbNF81OI?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/XSmBfn462wU?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/WYHeW73tA5s?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/D9UB4sSIWzw?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/FUXGg0gTmzY?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/TXZh1sqBDKU?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/BJVr0eMUTSU?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/jhoYzh--tVw?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/VscpAyJMd98?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/ekbkIImHctQ?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
			
				
	<div class="contentdiv">
		<div class="fyts-videoWrapper">
		
		<iframe id="ytplayer" width="100%" height="100%" src="https://www.youtube.com/embed/Y1jafS4NSJM
?theme=light&color=red&autohide=0&showinfo=1&autoplay=0" frameborder="0" allowfullscreen /></iframe>
		 
		</div>
	</div>
	</div>

<div id="paginate-fytslider380" class="paginationfytslide">
	<div style="text-align: center;" class="paginationfytslide-inner">
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/dYqQQ8k8ETs/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/rGrPbNF81OI/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/XSmBfn462wU/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/WYHeW73tA5s/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/D9UB4sSIWzw/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/FUXGg0gTmzY/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/TXZh1sqBDKU/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/BJVr0eMUTSU/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/jhoYzh--tVw/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/VscpAyJMd98/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/ekbkIImHctQ/default.jpg" width="22%" height="auto"></img>
		</a>
			<a href="#" class="toc">
			<img src="https://i3.ytimg.com/vi/Y1jafS4NSJM
/default.jpg" width="22%" height="auto"></img>
		</a>
		</div>
	<div style="text-align: right; font-size:8px; padding-right:3px; font-family:fantasy; color:#800000;"><a href="http://showlands.com" target="_blank" title="Video System by Featured YouTube Slider">YouTube Slider</a></div>
</div>
</div>
<script type="text/javascript">

featuredcontentslider.init({
	id: "fytslider380",  //id of main slider DIV
	contentsource: ["inline", ""],  
	toc: "markup",  //Valid values: "#increment", "markup", ["label1", "label2", etc]
	nextprev: ["Previous", "Next"],  //labels for "prev" and "next" links. Set to "" to hide.
	revealtype: "click", //Behavior of pagination links to reveal the slides: "click" or "mouseover"
	enablefade: [true, 0.2],  //[true/false, fadedegree]
	autorotate: [false, 3000],  //[true/false, pausetime]
	onChange: function(previndex, curindex){  //event handler fired whenever script changes slide
		//previndex holds index of last slide viewed b4 current (1=1st slide, 2nd=2nd etc)
		//curindex holds index of currently shown slide (1=1st slide, 2nd=2nd etc)
	}
})

</script></div>
		
          
          </div>
	
    
                </div>
            </div>
            <!-- /sidebar -->
             
                           
		</div>
        
                <div id="icecarousel"> 
            
<div style="border: 0px !important;">
<div id="djslider-loader383" class="djslider-loader djslider-loader-default" data-animation='{"auto":"1","transition":"easeInOutExpo","css3transition":"cubic-bezier(1.000, 0.000, 0.000, 1.000)","duration":400,"delay":3400}' data-djslider='{"id":"383","slider_type":"0","slide_size":250,"visible_slides":"5","direction":"left","show_buttons":"1","show_arrows":"1","preload":"800","css3":"1"}' tabindex="0">
    <div id="djslider383" class="djslider djslider-default" style="height: 240px; width: 1240px; max-width: 1240px !important;">
        <div id="slider-container383" class="slider-container">
        	<ul id="slider383" class="djslider-in">
          		          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/1.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/1.png" alt="1.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/2.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/2.png" alt="2.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/3.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/3.png" alt="3.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/4.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/4.png" alt="4.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/5.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/5.png" alt="5.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/6.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/6.png" alt="6.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/7.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/7.png" alt="7.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/8.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/8.png" alt="8.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/9.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/9.png" alt="9.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/10.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/10.png" alt="10.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                          			<li style="margin: 0 10px 0px 0 !important; height: 240px; width: 240px;">
          					            											<a class="image-link" data-title="" href="/images/image_gallery/ICECARRUSEL/11.png" target="_self">
															<img class="dj-image" src="/images/image_gallery/ICECARRUSEL/11.png" alt="11.png" style="width: 100%; height: auto;"/>
															</a>
																									
						
					</li>
                        	</ul>
        </div>
                <div id="navigation383" class="navigation-container" style="top: 16.6666666667%; margin: 0 0.806451612903%;">
        	        	<img id="prev383" class="prev-button showOnHover" src="/modules/mod_djimageslider/themes/default/images/prev.png" alt="Previous" tabindex="0" />
			<img id="next383" class="next-button showOnHover" src="/modules/mod_djimageslider/themes/default/images/next.png" alt="Next" tabindex="0" />
									<img id="play383" class="play-button showOnHover" src="/modules/mod_djimageslider/themes/default/images/play.png" alt="Play" tabindex="0" />
			<img id="pause383" class="pause-button showOnHover" src="/modules/mod_djimageslider/themes/default/images/pause.png" alt="Pause" tabindex="0" />
			        </div>
                    </div>
</div>
</div>
<div class="djslider-end" style="clear: both" tabindex="0"></div>           
        </div>   
                </div>   

    </section>
    <!-- / Content  --> 

      
	<footer id="footer" class="container">
		
		 
		<div id="copyright">
        	<div>
                <p class="copytext">
                    &copy; 2018 FDIM 
                </p>          
                <ul class="nav menu">
<li class="item-538"><a href="/info@fdim.org.sv" >info@fdim.org.sv</a></li><li class="item-536"><a href="#" >Services</a></li><li class="item-537"><a href="#" >Contact</a></li><li class="item-743"><a href="http://www.icetheme.com" target="_blank" >Designed by IceTheme</a></li></ul>

      		</div>
		</div>
   
	</footer>   
  
	    <div id="gotop" class="">
        <a href="#" class="scrollup">Go Top</a>
    </div>
      

        
	






</body>
</html>