


<!DOCTYPE html>

<html xmlns="http://www.w3.org/1999/xhtml">
<head><link rel="stylesheet" type="text/css" href="/DXR.axd?r=0_1747,1_50,1_53,1_51,1_16,0_1750-OVpNf&p=7de66f31" /><link rel="stylesheet" type="text/css" href="/DXR.axd?r=0_5900-OVpNf" /><link rel="stylesheet" type="text/css" href="/DXR.axd?r=0_4860,0_4864,0_1856-OVpNf&p=7de66f31" /><link rel="stylesheet" type="text/css" href="/DXR.axd?r=0_1859,0_974,0_978-OVpNf&p=7de66f31" /><link rel="stylesheet" type="text/css" href="/DXR.axd?r=0_1757,0_1760,1_17,0_3417,0_3421-OVpNf&p=7de66f31" /><meta name="robots" content="all" /><meta name="viewport" content="width=device-width, initial-scale=1.0" /><title>
	Empleos Públicos en El Salvador
</title><link rel="shortcut icon" href="Content/Images/favicon.ico" /><meta name="Keywords" content="empleos,el salvador,puestos,trabajo,gobierno,tecnica,plazas,elsalvador,ofertas,san salvador,secretaria tecnica,gobierno abierto" /><meta name="description" content="El Gobierno de la República de El Salvador busca estandarizar y propiciar una transparente y eficiente gestión de los procesos de dotación, selección y ascensos, donde el mérito, la idoneidad, la igualdad de oportunidades y la no discriminación sean los elementos fundamentales." /><link href="//fonts.googleapis.com/css?family=Montserrat" rel="stylesheet" type="text/css" /><link rel="stylesheet" href="https://cdnjs.cloudflare.com/ajax/libs/font-awesome/4.7.0/css/font-awesome.min.css" /><link rel="stylesheet" type="text/css" href="Content/Site.css" />
<script>
    (function (i, s, o, g, r, a, m) {
        i['GoogleAnalyticsObject'] = r; i[r] = i[r] || function () {
            (i[r].q = i[r].q || []).push(arguments)
        }, i[r].l = 1 * new Date(); a = s.createElement(o),
        m = s.getElementsByTagName(o)[0]; a.async = 1; a.src = g; m.parentNode.insertBefore(a, m)
    })(window, document, 'script', 'https://www.google-analytics.com/analytics.js', 'ga');

    ga('create', 'UA-71404431-1', 'auto');
    ga('send', 'pageview');

</script>
</head>
<body>
   <form method="post" action="./" id="aspnetForm">
<input type="hidden" name="__VIEWSTATE" id="__VIEWSTATE" value="/wEPDwUKMjEwMzgwMTg1OA9kFgJmD2QWAgIDD2QWCAIBD2QWAgIBD2QWAgIBDzwrAAoBAA8WAh4OXyFVc2VWaWV3U3RhdGVnZGQCAw9kFgJmDzwrAAoCAA8WAh8AZ2QGD2QQFgFmFgE8KwAMAQAWAh4IU2VsZWN0ZWRnZGQCBQ9kFhICAQ8WAh4EVGV4dAUBMGQCAw8WAh8CBQEwZAIFDxYCHwIFATJkAgcPFgIfAgUBNmQCCw8WAh8CBQUxLDM4OGQCDQ8WAh8CBQ8yNiBWYWNhbnRlcyBlbiBkAg8PFgIfAgUCMjZkAhEPFgIfAgUKMTUsOTc0LDgwNmQCEw9kFgQCAQ88KwAIAQAPFgIfAGdkZAIDDzwrACYDAA8WAh4PRGF0YVNvdXJjZUJvdW5kZ2QGD2QQFgdmAgECAgIDAgQCBQIGFgc8KwAMAQAWAh4LR2xvYmFsSW5kZXhmPCsADAEAFgIfBAIBPCsADAEAFgIfBAICPCsADAEAFgIfBAIDPCsADAEAFgIfBAIEPCsADAEAFgIfBAIFPCsADAEAFgIfBAIGDxYHAgECAQIBAgECAQIBAgEWAQV/RGV2RXhwcmVzcy5XZWIuR3JpZFZpZXdEYXRhVGV4dENvbHVtbiwgRGV2RXhwcmVzcy5XZWIudjE3LjIsIFZlcnNpb249MTcuMi4zLjAsIEN1bHR1cmU9bmV1dHJhbCwgUHVibGljS2V5VG9rZW49Yjg4ZDE3NTRkNzAwZTQ5YRg8KwAHAQUUKwACZGQWAgIBD2QWAmYPZBYCZg9kFgJmD2QWAgULRFhNYWluVGFibGUPZBYKBQpEWERhdGFSb3cwD2QWAgUJdGNjZWxsMF8wD2QWAmYPZBYCZg9kFgJmDxUCBDE5MjUqQXNpc3RlbnRlIGRlIEdlc3Rpw7NuIERvY3VtZW50YWwgeSBBcmNoaXZvZAUKRFhEYXRhUm93MQ9kFgIFCXRjY2VsbDFfMA9kFgJmD2QWAmYPZBYCZg8VAgQyMDYxEVBvcnRlcm8gVmlnaWxhbnRlZAUKRFhEYXRhUm93Mg9kFgIFCXRjY2VsbDJfMA9kFgJmD2QWAmYPZBYCZg8VAgQyMDYyFEF1eGlsaWFyIGRlIFNlcnZpY2lvZAUKRFhEYXRhUm93Mw9kFgIFCXRjY2VsbDNfMA9kFgJmD2QWAmYPZBYCZg8VAgQyMDYwDE1vdG9yaXN0YSBJSWQFCkRYRGF0YVJvdzQPZBYCBQl0Y2NlbGw0XzAPZBYCZg9kFgJmD2QWAmYPFQIEMjA1OQxNb3RvcmlzdGEgSUlkAgcPPCsACQEADxYCHwBnZGQYAgUeX19Db250cm9sc1JlcXVpcmVQb3N0QmFja0tleV9fFhUFFmN0bDAwJGJ0bklkZW50aWZpY2Fyc2UFF2N0bDAwJHVjTWVudSRIZWFkZXJNZW51BR1jdGwwMCRNYWluQ29udGVudCRBU1B4QnV0dG9uMQUuY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkcGFuZWxJbnMkMzEwOAUuY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkcGFuZWxJbnMkNDIwMwUuY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkcGFuZWxJbnMkMDcwMgUuY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkcGFuZWxJbnMkMjMwMwUsY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkcGFuZWxJbnMkMzIFNmN0bDAwJE1haW5Db250ZW50JHVsdGltb3NFbXBsZW9zJGdyaWRQdWVzdG9zUHVibGljYWRvcwVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwwXzUkYnRuQXBsaWNhcgVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwwXzUkYnRuUHJvY2VzbwVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwxXzUkYnRuQXBsaWNhcgVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwxXzUkYnRuUHJvY2VzbwVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwyXzUkYnRuQXBsaWNhcgVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwyXzUkYnRuUHJvY2VzbwVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwzXzUkYnRuQXBsaWNhcgVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGwzXzUkYnRuUHJvY2VzbwVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGw0XzUkYnRuQXBsaWNhcgVJY3RsMDAkTWFpbkNvbnRlbnQkdWx0aW1vc0VtcGxlb3MkZ3JpZFB1ZXN0b3NQdWJsaWNhZG9zJGNlbGw0XzUkYnRuUHJvY2VzbwUSY3RsMDAkcG9wdXBNZW5zYWplBR9jdGwwMCRwb3B1cE1lbnNhamUkVFBDRm0xJGJ0bk9rBRBjdGwwMCRNdWx0aVZpZXcxDw9kZmR4YBLI2FUxRfo+YMLdZSmbjIqBDW53UO1B0qQwBtYOqQ==" />

<input type="hidden" name="__VIEWSTATEGENERATOR" id="__VIEWSTATEGENERATOR" value="CA0B0334" />
<input type="hidden" name="__PREVIOUSPAGE" id="__PREVIOUSPAGE" value="VUkEeIPvU_tHiE7oCIu6Q9dEAx9EBR9QmJXr25KT4deU-aayE7-aWfId-jeqiNv2I9JMsj2Jgn5Z80c-Bj5ZMkGQVVwUmsPaBMqmzO8qkVc1" />
<input type="hidden" name="__EVENTVALIDATION" id="__EVENTVALIDATION" value="/wEdAAORNVbo5RxNLY70PEqYcrmDx9IsQjaMxk+v7T5d+FERI2zc5M1SDvhoZPdfj1GZlzMCiib+aluH5MJ4K0SiRM/HhPHfhUnfQP++sx71qw9GZg==" />
   <div id="inicio">
    <div id="top">
        <div id="top-container">
            <div id="logo" class="top-item"></div>
            <div id="titulo" class="top-item">Empleos Públicos en El Salvador</div>
            <div id="login" class="top-item">
                

                            <input type="hidden"/><script id="dxis_929767809" src="/DXR.axd?r=1_304,1_185,1_298,1_211,1_221,1_188,1_182,1_198,1_290,1_296,1_279,1_196,1_254,1_256,1_263,1_235,1_248,1_244,1_242,1_251,1_238,1_239,1_247,1_209,1_217,1_224,1_288-MVpNf" type="text/javascript"></script><div title="Identificación si ya se tiene usuario y clave" class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_btnIdentificarse" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
	<div class="dxb">
		<input id="ctl00_btnIdentificarse_I" title="Identificación si ya se tiene usuario y clave" class="dxb-hb" value="Iniciar Sesión" type="button" name="ctl00$btnIdentificarse" /><img class="dx-vam" src="Content/Images/Employee_16x16.png" alt="" style="margin-right:4px;" /><span class="dx-vam">Iniciar Sesi&#243;n</span>
	</div>
</div><script id="dxss_1611404372" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_btnIdentificarse',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_btnIdentificarse',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_btnIdentificarse',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_btnIdentificarse','',{'autoPostBack':true,'uniqueID':'ctl00$btnIdentificarse','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$btnIdentificarse",  postBackArg, true, "", "Login.aspx", false, true)); }});

//-->
</script>
                    
            </div>
        </div>
        <div id="top-menu">
            <div class="dxmLite_PlasticBlue dxm-ltr">
	<div class="dxm-main dxm-horizontal dxm-noWrap headerMenu" id="ctl00_ucMenu_HeaderMenu" style="border-top-width:1px;padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;">
		<ul class="dx dxm-image-l">
			<li class="dxm-item dxm-selected dxm-noSubMenu"><div class="dxm-content dxm-hasText">
				<img class="dxm-image dx-vam" src="Content/Images/Home_32x32.png" alt="" /><span class="dx-vam">Inicio</span>
			</div></li><li class="dxm-separator"><b></b></li><li class="dxm-item dxm-noSubMenu"><a class="dxm-content dxm-hasText dx" href="Concursos.aspx"><img class="dxm-image dx-vam" src="Content/Images/Concurso.png" alt="" /><span class="dx-vam">Concursos</span></a></li><li class="dxm-separator"><b></b></li><li class="dxm-item dxm-noSubMenu"><a class="dxm-content dxm-hasText dx" href="Registro.aspx"><img class="dxm-image dx-vam" src="Content/Images/Menu.png" alt="" /><span class="dx-vam">Registrate</span></a></li><li class="dxm-separator"><b></b></li><li class="dxm-item dxm-noSubMenu"><a class="dxm-content dxm-hasText dx" href="wfEstadistica.aspx"><img class="dxm-image dx-vam" src="Content/Images/Chart2_32x32.png" alt="" /><span class="dx-vam">Estad&#237;sticas</span></a></li><li class="dxm-separator"><b></b></li><li class="dxm-item dxm-noSubMenu"><a class="dxm-content dxm-hasText dx" href="wfContacto.aspx"><img class="dxm-image dx-vam" src="Content/Images/Question.png" alt="" /><span class="dx-vam">Soporte</span></a></li><li class="dxm-spacing dxm-amis"></li><li class="dxm-item dxm-dropDownMode dxm-noImage dxm-ami"><div class="dxm-content" style="padding-right:13px;">
				<span class="dx-vam">&nbsp;</span>
			</div><div class="dxm-popOut">
				<img class="dxWeb_mAdaptiveMenu_PlasticBlue dxm-pImage" src="/DXR.axd?r=1_58-MVpNf" alt="..." />
			</div></li>
		</ul>
	</div><b class="dx-clear"></b><div id="ctl00_ucMenu_HeaderMenu_DXM5_" style="z-index:20000;display:none;">
		<div class="dxm-shadow dxm-popup dxm-am">
			<ul class="dx dxm-gutter">

			</ul>
		</div>
	</div>
</div><script id="dxss_1961056024" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_ucMenu_HeaderMenu',[[[''],[''],['DXI0_'],['','T']],[['dxm-hovered',''],['',''],['DXI1_','DXI2_','DXI3_','DXI4_'],['','T']],[['dxm-hovered','',''],['','',''],['DXI5_'],['','P','T']],[[''],[''],['DXME5_','DXMBC5_']]]);
ASPx.AddDisabledItems('ctl00_ucMenu_HeaderMenu',[[['dxm-disabled'],[''],['DXI0_','DXI1_','DXI2_','DXI3_','DXI4_'],['','T']],[['dxm-disabled'],[''],['DXI5_'],['','P','T']]]);
ASPx.createControl(ASPxClientMenu,'ctl00_ucMenu_HeaderMenu','headerMenu',{'uniqueID':'ctl00$ucMenu$HeaderMenu','renderData':{'':[0,[1],[2],[3],[4],5]},'subMenuFIYOffset':-1,'subMenuLIYOffset':-1,'subMenuYOffset':-1,'rootSubMenuFIXOffset':1,'rootSubMenuLIXOffset':1,'rootSubMenuXOffset':1},null,null,{'items':[{},{},{},{},{},{}],'adaptiveModeData':5});

//-->
</script>
        </div>
    </div>
                    
    <div id="banner">
        <div id="tableBanner">
                    <div class="flex-contador">
                        <span class="label">0</span>
                        <span class="label">0</span>
                        <span class="label">2</span>
                        <span class="label">6</span>
                    </div>

                <div class="bannerTitulo">Empleos públicos disponibles</div>
                    <div class="bannerSubTitulo">El Gobierno de la República de El Salvador busca estandarizar y propiciar una transparente y eficiente gestión de los procesos de dotación, selección y ascensos, donde el mérito, la idoneidad, la igualdad de oportunidades y la no discriminación sean los elementos fundamentales.</div>
                    <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ASPxButton1" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
	<div class="dxb">
		<input id="ctl00_MainContent_ASPxButton1_I" class="dxb-hb" value="Consultar Listado de Concursos" type="button" name="ctl00$MainContent$ASPxButton1" /><span class="dx-vam">Consultar Listado de Concursos</span>
	</div>
</div><script id="dxss_844865710" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ASPxButton1',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ASPxButton1',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ASPxButton1',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ASPxButton1',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ASPxButton1','',{'uniqueID':'ctl00$MainContent$ASPxButton1','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ASPxButton1",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {
	window.location = "Concursos.aspx";
}});

//-->
</script>

                <div class="flex-container">
                    <div class="flex-item">
                          <img src="Content/Images/maletin.png" />
                            <div class="bannerText">
                                1,388
                                <br />Concursos a la fecha
                            </div>
                    </div>
                    <div class="flex-item">
                        <img src="Content/Images/icon-sales.png" />
                        <div class="bannerText">
                                26 Vacantes en <br />26 Concursos disponibles
                            </div>
                    </div>
                    <div class="flex-item">
                       <img src="Content/Images/icon-statistics.png" />
                        <div class="bannerText">
                                15,974,806<br />Visitas a la fecha
                            </div>
                    </div>
                </div>

            
        </div>

        
    </div>
    <div id="content">
        <div id="content-wrap">
    
<script type="text/javascript">
     // <![CDATA[
        function OnMoreInfoClick(key) {
            
            window.location.href = 'wfPlaza.aspx?p=' + key;
        }
        function Proceso(key) {

            window.location.href = 'wfProceso.aspx?p=' + key;
        }

     function CallForm(key) {
         popupPlaza.Show();
         cbpPlaza.PerformCallback(key);
     }
     // ]]> 
</script>
<table style="width:100%">
    <tr>
        <td style="width:20%;vertical-align:top;" class="lateral">
            <h3 style="text-align:left">Instituciones</h3>
            <div class="dxpnlControl_MaterialCompact" id="ctl00_MainContent_ultimosEmpleos_panelIns">
	<div title="Consejo Nacional de la Niñez y de la Adolescencia" class="dxbButton_Glass dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_panelIns_3108" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
		<div class="dxb">
			<input id="ctl00_MainContent_ultimosEmpleos_panelIns_3108_I" title="Consejo Nacional de la Niñez y de la Adolescencia" class="dxb-hb" value="CONNA" type="button" name="ctl00$MainContent$ultimosEmpleos$panelIns$3108" /><span class="dx-vam">CONNA</span>
		</div>
	</div><script id="dxss_724830862" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_panelIns_3108',[[['dxbButtonHover_Glass'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_panelIns_3108',[[['dxbButtonPressed_Glass'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_panelIns_3108',[[['dxbDisabled_Glass'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_panelIns_3108',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_panelIns_3108','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$panelIns$3108','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$panelIns$3108",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e)  { window.location = 'Concursos.aspx?ins=3108'; }});

//-->
</script><div title="Escuela Nacional de Agricultura" class="dxbButton_Glass dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_panelIns_4203" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
		<div class="dxb">
			<input id="ctl00_MainContent_ultimosEmpleos_panelIns_4203_I" title="Escuela Nacional de Agricultura" class="dxb-hb" value="ENA" type="button" name="ctl00$MainContent$ultimosEmpleos$panelIns$4203" /><span class="dx-vam">ENA</span>
		</div>
	</div><script id="dxss_1689557998" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_panelIns_4203',[[['dxbButtonHover_Glass'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_panelIns_4203',[[['dxbButtonPressed_Glass'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_panelIns_4203',[[['dxbDisabled_Glass'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_panelIns_4203',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_panelIns_4203','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$panelIns$4203','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$panelIns$4203",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e)  { window.location = 'Concursos.aspx?ins=4203'; }});

//-->
</script><div title="Instituto Nacional de Pensiones de los Empleados Públicos" class="dxbButton_Glass dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_panelIns_0702" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
		<div class="dxb">
			<input id="ctl00_MainContent_ultimosEmpleos_panelIns_0702_I" title="Instituto Nacional de Pensiones de los Empleados Públicos" class="dxb-hb" value="INPEP" type="button" name="ctl00$MainContent$ultimosEmpleos$panelIns$0702" /><span class="dx-vam">INPEP</span>
		</div>
	</div><script id="dxss_2033176814" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_panelIns_0702',[[['dxbButtonHover_Glass'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_panelIns_0702',[[['dxbButtonPressed_Glass'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_panelIns_0702',[[['dxbDisabled_Glass'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_panelIns_0702',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_panelIns_0702','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$panelIns$0702','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$panelIns$0702",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e)  { window.location = 'Concursos.aspx?ins=0702'; }});

//-->
</script><div title="Instituto Salvadoreño de Desarrollo Municipal" class="dxbButton_Glass dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_panelIns_2303" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
		<div class="dxb">
			<input id="ctl00_MainContent_ultimosEmpleos_panelIns_2303_I" title="Instituto Salvadoreño de Desarrollo Municipal" class="dxb-hb" value="ISDEM" type="button" name="ctl00$MainContent$ultimosEmpleos$panelIns$2303" /><span class="dx-vam">ISDEM</span>
		</div>
	</div><script id="dxss_2123822898" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_panelIns_2303',[[['dxbButtonHover_Glass'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_panelIns_2303',[[['dxbButtonPressed_Glass'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_panelIns_2303',[[['dxbDisabled_Glass'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_panelIns_2303',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_panelIns_2303','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$panelIns$2303','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$panelIns$2303",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e)  { window.location = 'Concursos.aspx?ins=2303'; }});

//-->
</script><div title="Ministerio de Salud" class="dxbButton_Glass dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_panelIns_32" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
		<div class="dxb">
			<input id="ctl00_MainContent_ultimosEmpleos_panelIns_32_I" title="Ministerio de Salud" class="dxb-hb" value="MINSAL" type="button" name="ctl00$MainContent$ultimosEmpleos$panelIns$32" /><span class="dx-vam">MINSAL</span>
		</div>
	</div><script id="dxss_1478111154" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_panelIns_32',[[['dxbButtonHover_Glass'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_panelIns_32',[[['dxbButtonPressed_Glass'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_panelIns_32',[[['dxbDisabled_Glass'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_panelIns_32',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_panelIns_32','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$panelIns$32','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$panelIns$32",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e)  { window.location = 'Concursos.aspx?ins=32'; }});

//-->
</script>
</div>
        </td>
        <td style="width:80%;padding-left:10px;vertical-align:top;">
            <h3 style="text-align:left">Últimos concursos publicados:</h3>
            <table class="dxgvControl_MaterialCompact dxgv" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados" width="100%" style="border-collapse:separate;">
	<tr>
		<td style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><div id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAHeaderPanel" class="dxgvAdaptiveHeaderPanel_MaterialCompact" oncontextmenu="return ASPx.GVContextMenu(&#39;ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados&#39;,event);" style="display:none;">
			<div id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXADHeader" class="dxgvADH" style="display:none;">
				<table>
					<tr class="dxgvADHTR">
						<td></td>
					</tr>
				</table>
			</div>
		</div><table id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXMainTable" class="dxgvTable_MaterialCompact" onclick="ASPx.GTableClick(&#39;ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados&#39;, event);" ondblclick="ASPx.GVTableDblClick(&#39;ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados&#39;, event);" oncontextmenu="return ASPx.GVContextMenu(&#39;ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados&#39;,event);" width="100%" style="empty-cells:show;">
			<tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXHeadersRow0">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col0" title="Nombre del puesto funcional en el Gobierno" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="33%" style="border-top-width:0px;border-left-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap">Título del Puesto</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col1" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="10%" style="border-top-width:0px;border-left-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap">Institución</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col3" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="5%" style="text-align:Center;border-top-width:0px;border-left-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap" style="text-align:Center;">Salario</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col2" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="7%" style="border-top-width:0px;border-left-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap">Vacantes</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col4" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="15%" style="text-align:Center;border-top-width:0px;border-left-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap" style="text-align:Center;">Ubicación</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_col5" class="dxgvHeader_MaterialCompact hide-header dx-wrap" width="30%" style="text-align:Center;border-top-width:0px;border-left-width:0px;border-right-width:0px;cursor:default;"><table width="100%">
					<tr>
						<td class="dx-wrap" style="text-align:Center;">Acción</td><td width="1" style="text-align:right;"><span class="dx-vam">&nbsp;</span></td>
					</tr>
				</table></td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXADRow" class="dxgvDetailRow_MaterialCompact dxgvADR" style="display:none;">
				<td class="dxgv dxgvDetailCell_MaterialCompact" colspan="6"><div class="dxflFormLayout_MaterialCompact dxflViewFormLayoutSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL">
					<table class="dxflGroup_MaterialCompact dxflGroupSys dxflAGSys" style="border-collapse:separate;">
						<tr>
							<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_0" class="dxflGroupCell_MaterialCompact" colspan="2" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><table class="dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact" style="border-collapse:separate;">
								<tr>
									<td class="dxflHALSys dxflVATSys dxflCaptionCell_MaterialCompact dxflCaptionCellSys dxgvADCC"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_0_Cap" class="dxDefaultCursor dxflCaption_MaterialCompact">T&#237;tulo del Puesto:</span></td>
								</tr><tr>
									<td class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC0">&nbsp;</td>
								</tr>
							</table></td>
						</tr><tr>
							<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_1" class="dxflGroupCell_MaterialCompact" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><table class="dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact" style="border-collapse:separate;">
								<tr>
									<td class="dxflHALSys dxflVATSys dxflCaptionCell_MaterialCompact dxflCaptionCellSys dxgvADCC"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_1_Cap" class="dxDefaultCursor dxflCaption_MaterialCompact">Instituci&#243;n:</span></td>
								</tr><tr>
									<td class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC1">&nbsp;</td>
								</tr>
							</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_2" class="dxflGroupCell_MaterialCompact" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><table class="dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact" style="border-collapse:separate;">
								<tr>
									<td class="dxflHALSys dxflVATSys dxflCaptionCell_MaterialCompact dxflCaptionCellSys dxgvADCC"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_2_Cap" class="dxDefaultCursor dxflCaption_MaterialCompact">Salario:</span></td>
								</tr><tr>
									<td class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC3">&nbsp;</td>
								</tr>
							</table></td>
						</tr><tr>
							<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_3" class="dxflGroupCell_MaterialCompact" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><table class="dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact" style="border-collapse:separate;">
								<tr>
									<td class="dxflHALSys dxflVATSys dxflCaptionCell_MaterialCompact dxflCaptionCellSys dxgvADCC"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_3_Cap" class="dxDefaultCursor dxflCaption_MaterialCompact">Vacantes:</span></td>
								</tr><tr>
									<td class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC2">&nbsp;</td>
								</tr>
							</table></td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_4" class="dxflGroupCell_MaterialCompact" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><table class="dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact" style="border-collapse:separate;">
								<tr>
									<td class="dxflHALSys dxflVATSys dxflCaptionCell_MaterialCompact dxflCaptionCellSys dxgvADCC"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_4_Cap" class="dxDefaultCursor dxflCaption_MaterialCompact">Ubicaci&#243;n:</span></td>
								</tr><tr>
									<td class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC4">&nbsp;</td>
								</tr>
							</table></td>
						</tr><tr>
							<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL_5" class="dxflGroupCell_MaterialCompact" colspan="2" style="padding-left:0px;padding-right:0px;padding-top:0px;padding-bottom:0px;"><div class="dxflNestedControlCell_MaterialCompact dxgvADDC dxgvADLIC5 dxflCLTSys dxflItemSys dxflTextItemSys dxflItem_MaterialCompact">
								&nbsp;
							</div></td>
						</tr>
					</table>
				</div><script id="dxss_1152669692" type="text/javascript">
<!--
ASPx.createControl(ASPxClientFormLayout,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXAFL','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$DXAFL'});

//-->
</script></td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXDataRow0" class="dxgvDataRow_MaterialCompact">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell0_0" class="dxgv">
                    <a href="javascript:void(0);" onclick="OnMoreInfoClick('1925')" class="mayusculas">
                        Asistente de Gestión Documental y Archivo
                    </a>
                </td><td title="Instituto Salvadoreño de Desarrollo Municipal" class="dxgv">ISDEM</td><td class="dxgv dx-ar">$400.00</td><td class="dxgv dx-ar">1</td><td class="dxgv dx-ac">SAN SALVADOR</td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell0_5" class="dxgv dx-ac" style="border-right-width:0px;">
                                <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar_I" class="dxb-hb" value="Aplicar" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnAplicar" /><span class="dx-vam">Aplicar</span>
					</div>
				</div><script id="dxss_1822974127" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnAplicar','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnAplicar','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnAplicar",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {OnMoreInfoClick('1925');}});

//-->
</script>
                                <div class="dxbButton_Office2003Silver dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso_I" class="dxb-hb" value="Ver proceso" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnProceso" /><span class="dx-vam">Ver proceso</span>
					</div>
				</div><script id="dxss_1645733831" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso',[[['dxbButtonHover_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso',[[['dxbButtonPressed_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso',[[['dxbDisabled_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell0_5_btnProceso','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnProceso','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell0_5$btnProceso",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {Proceso('1925');}});

//-->
</script>
                </td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXDataRow1" class="dxgvDataRow_MaterialCompact dxgvDataRowAlt_MaterialCompact">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell1_0" class="dxgv">
                    <a href="javascript:void(0);" onclick="OnMoreInfoClick('2061')" class="mayusculas">
                        Portero Vigilante
                    </a>
                </td><td title="Ministerio de Salud" class="dxgv">MINSAL</td><td class="dxgv dx-ar">$286.29</td><td class="dxgv dx-ar">1</td><td class="dxgv dx-ac">SAN VICENTE</td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell1_5" class="dxgv dx-ac" style="border-right-width:0px;">
                                <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar_I" class="dxb-hb" value="Aplicar" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnAplicar" /><span class="dx-vam">Aplicar</span>
					</div>
				</div><script id="dxss_1076012822" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnAplicar','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnAplicar','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnAplicar",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {OnMoreInfoClick('2061');}});

//-->
</script>
                                <div class="dxbButton_Office2003Silver dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso_I" class="dxb-hb" value="Ver proceso" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnProceso" /><span class="dx-vam">Ver proceso</span>
					</div>
				</div><script id="dxss_1814137480" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso',[[['dxbButtonHover_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso',[[['dxbButtonPressed_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso',[[['dxbDisabled_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell1_5_btnProceso','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnProceso','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell1_5$btnProceso",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {Proceso('2061');}});

//-->
</script>
                </td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXDataRow2" class="dxgvDataRow_MaterialCompact">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell2_0" class="dxgv">
                    <a href="javascript:void(0);" onclick="OnMoreInfoClick('2062')" class="mayusculas">
                        Auxiliar de Servicio
                    </a>
                </td><td title="Ministerio de Salud" class="dxgv">MINSAL</td><td class="dxgv dx-ar">$256.58</td><td class="dxgv dx-ar">1</td><td class="dxgv dx-ac">SAN ISIDRO</td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell2_5" class="dxgv dx-ac" style="border-right-width:0px;">
                                <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar_I" class="dxb-hb" value="Aplicar" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnAplicar" /><span class="dx-vam">Aplicar</span>
					</div>
				</div><script id="dxss_1458568100" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnAplicar','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnAplicar','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnAplicar",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {OnMoreInfoClick('2062');}});

//-->
</script>
                                <div class="dxbButton_Office2003Silver dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso_I" class="dxb-hb" value="Ver proceso" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnProceso" /><span class="dx-vam">Ver proceso</span>
					</div>
				</div><script id="dxss_1505674914" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso',[[['dxbButtonHover_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso',[[['dxbButtonPressed_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso',[[['dxbDisabled_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell2_5_btnProceso','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnProceso','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell2_5$btnProceso",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {Proceso('2062');}});

//-->
</script>
                </td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXDataRow3" class="dxgvDataRow_MaterialCompact dxgvDataRowAlt_MaterialCompact">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell3_0" class="dxgv">
                    <a href="javascript:void(0);" onclick="OnMoreInfoClick('2060')" class="mayusculas">
                        Motorista II
                    </a>
                </td><td title="Ministerio de Salud" class="dxgv">MINSAL</td><td class="dxgv dx-ar">$292.58</td><td class="dxgv dx-ar">1</td><td class="dxgv dx-ac">SAN VICENTE</td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell3_5" class="dxgv dx-ac" style="border-right-width:0px;">
                                <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar_I" class="dxb-hb" value="Aplicar" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnAplicar" /><span class="dx-vam">Aplicar</span>
					</div>
				</div><script id="dxss_498767943" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnAplicar','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnAplicar','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnAplicar",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {OnMoreInfoClick('2060');}});

//-->
</script>
                                <div class="dxbButton_Office2003Silver dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso_I" class="dxb-hb" value="Ver proceso" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnProceso" /><span class="dx-vam">Ver proceso</span>
					</div>
				</div><script id="dxss_1333176385" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso',[[['dxbButtonHover_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso',[[['dxbButtonPressed_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso',[[['dxbDisabled_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell3_5_btnProceso','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnProceso','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell3_5$btnProceso",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {Proceso('2060');}});

//-->
</script>
                </td>
			</tr><tr id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_DXDataRow4" class="dxgvDataRow_MaterialCompact">
				<td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell4_0" class="dxgv" style="border-bottom-width:0px;">
                    <a href="javascript:void(0);" onclick="OnMoreInfoClick('2059')" class="mayusculas">
                        Motorista II
                    </a>
                </td><td title="Ministerio de Salud" class="dxgv" style="border-bottom-width:0px;">MINSAL</td><td class="dxgv dx-ar" style="border-bottom-width:0px;">$292.58</td><td class="dxgv dx-ar" style="border-bottom-width:0px;">1</td><td class="dxgv dx-ac" style="border-bottom-width:0px;">SAN VICENTE</td><td id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_tccell4_5" class="dxgv dx-ac" style="border-right-width:0px;border-bottom-width:0px;">
                                <div class="dxbButton_MaterialCompact dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar_I" class="dxb-hb" value="Aplicar" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnAplicar" /><span class="dx-vam">Aplicar</span>
					</div>
				</div><script id="dxss_1434691368" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnAplicar','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnAplicar','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnAplicar",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {OnMoreInfoClick('2059');}});

//-->
</script>
                                <div class="dxbButton_Office2003Silver dxbButtonSys dxbTSys" id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
					<div class="dxb">
						<input id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso_I" class="dxb-hb" value="Ver proceso" type="button" name="ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnProceso" /><span class="dx-vam">Ver proceso</span>
					</div>
				</div><script id="dxss_1084600010" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso',[[['dxbButtonHover_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso',[[['dxbButtonPressed_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso',[[['dxbDisabled_Office2003Silver'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_cell4_5_btnProceso','',{'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnProceso','useSubmitBehavior':false,'autoPostBackFunction':function(postBackArg) { WebForm_DoPostBackWithOptions(new WebForm_PostBackOptions("ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados$cell4_5$btnProceso",  postBackArg, true, "", "", false, true)); }},{'Click':function(s, e) {Proceso('2059');}});

//-->
</script>
                </td>
			</tr>
		</table><table id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_LP" class="dxgvLoadingPanel_MaterialCompact" style="left:0px;top:0px;z-index:30000;display:none;">
			<tr>
				<td class="dx" style="padding-right:0px;"><img class="dxlp-loadingImage dxlp-imgPosLeft" src="/DXR.axd?r=1_58-MVpNf" alt="" style="vertical-align:middle;" /></td><td class="dx" style="padding-left:0px;"><span id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_TL">Cargando&hellip;</span></td>
			</tr>
		</table><div id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_LD" class="dxgvLoadingDiv_MaterialCompact" style="display:none;z-index:29999;position:absolute;">

		</div><img id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_IADD" class="dxGridView_gvDragAndDropArrowDown_MaterialCompact" src="/DXR.axd?r=1_58-MVpNf" alt="|" style="position:absolute;visibility:hidden;top:-100px;" /><img id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_IADU" class="dxGridView_gvDragAndDropArrowUp_MaterialCompact" src="/DXR.axd?r=1_58-MVpNf" alt="|" style="position:absolute;visibility:hidden;top:-100px;" /><img id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_IADL" class="dxGridView_gvDragAndDropArrowLeft_MaterialCompact" src="/DXR.axd?r=1_58-MVpNf" alt="|" style="position:absolute;visibility:hidden;top:-100px;" /><img id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_IADR" class="dxGridView_gvDragAndDropArrowRight_MaterialCompact" src="/DXR.axd?r=1_58-MVpNf" alt="|" style="position:absolute;visibility:hidden;top:-100px;" /><img id="ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados_IDHF" class="dxGridView_gvDragAndDropHideColumn_MaterialCompact" src="/DXR.axd?r=1_58-MVpNf" alt="Ocultar" style="position:absolute;visibility:hidden;top:-100px;" /></td>
	</tr>
</table><script id="dxss_2012138090" type="text/javascript">
<!--
ASPx.createControl(ASPxClientGridView,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados','gridPuestosPublicados',{'callBack':function(arg) { WebForm_DoCallback('ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados',arg,ASPx.Callback,'ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados',ASPx.CallbackError,true); },'uniqueID':'ctl00$MainContent$ultimosEmpleos$gridPuestosPublicados','stateObject':{'keys':['1925','2061','2062','2060','2059'],'callbackState':'qsnz0Wtk7HJZlCmMRmrc/g05mZhnbVnqZdXZgjOEsPs3YtGUg8J1aajI4/CmIPJpeDXAVXoQkf0CUOdUrkIkFC2Qxml7+l2l+LO9XiGQqq4Hcyy6d6DajxYzQiyWdILPtGGy0h09E0ogDLYbNopnQK37Bw+YTyFCyKNLiGVafYA2wODDt9irDA7So1r4zLvJFVoVnBYwqdllvkJRbE9EB+Qdwrg//Td7CAIX3oFBzZrUtfZOv+ql4hHvDwSWXJsLEROG7SVnDbhUVpmL0IA11aHXsydNd76rm32dVfw0bxdJgxof5o4hQX46cE9EIFAwK/ZhyC8FMLnCs7RsFcmI+9L+jIZoo+zsLSp5wl3Z/Vb7QjQgu/esT+/g6HGNaAOcHsNCSHumWTEB8v8QgITa+ynsgh1MrztVywlPFFfUUxcmiJkkz08oznGr3C5WaH4ut96f+usQclnL2YGie3KGwRk/wgV8dzmkBNYJIfVDAOuD/5El04v4IGQw8qGpDK/wXQByvJPtXAILqf0Lfxuehz84orri8m3C7gxn9JSNZ69utel+sB26ycHt1nSnMjNoKtrBv4DW5eyDbcqg9VWkz3qx0mWGEc3h1eJHgBhEqdc+PsxeC2wVd3qcXgCrz/hnUkaUK7O1YuZXJgMpNC3gjLBLz9TxJtCtIk7cG7w2LNvcAq7UH1bFd8HnHGHOcalkJcOgqbpuUB3WU1DEjyhodXaRhSbTKjfoeDxxqVX9DaVyQubxPgqSG69SNwwRWUx8L44avn8KukGvUNQohk20Xw2VLsdqMgVSL3oLJp+usClayNFwd7wk+eC8Wsj8ofujiieWSnxjYvq1PUcOPfmIrV00PC5ZJFphC8YKJfSCTZL7tSMhFtVQQmxS1WB0K2atmwocCEZN0SxybbLGJBvhzEnmHl+4mRyP490xbmopzimdcIvRd8HI1VZcAkTKwZNZQUhe8oqm9oGa1Qy/ZcZiAmOUUtxp9bJEPHjrdoZI4P65lPnnGaidNellwnyrHZm/fe1lWGPUuyoIxLM9ecyfu2nXyxAVKzVtprXr9vZUSURMOXS1BzM53HuIsVsEMedU1b/PSXJ18uKlUBSoZAHxtxXvRKPH6b+TxaLFK12X2DMnqGj1snXVkeDMjg4oWMzpJIeb0QpuJpLgItkrp2np6424075izyG67CDFYjGHqXHBk9cdUErEZmfMEKGH7YkcOd12ocFI5D18pprxwYlfFJ0ZSIktmcOrfmmDAYG8N9kcOV3cycxvTAhOnn+CJ8LAQpTpNMRg/0eKvvminNC1xxCff8prJFayG4hhaYyENrohflQHxbFJyct8opBSbGsJ379ijCN67syFCLPyGMjoH+8MAIDvBns6K6MvJVVqbSIqDHYCJYuTmddjy/YmR/P4NV7DB9tP5OMfJTcPddcpozPotWsY4CyhUUfNw9dtjL4MhP7sklNrU2Hd4kimMxDldooX/WLHmn7eEn/od87A9S73qJR9mFDDGE0yxu0P+EuJ57F2E4hpwFoQAVpqGDrHsXRXk/M2NQKCqcyIMPfG4LSmJF6ifxz2jK9D9TJczws7ocaKYrWDgFtkhADdfBBUCLGjqipvtY5GPtoJktZW+g==','selection':''},'callBacksEnabled':true,'pageRowCount':5,'pageRowSize':10,'pageIndex':-1,'pageCount':1,'selectedWithoutPageRowCount':0,'visibleStartIndex':0,'focusedRowIndex':-1,'allowFocusedRow':false,'allowSelectByItemClick':false,'allowSelectSingleRowOnly':false,'callbackOnFocusedRowChanged':false,'callbackOnSelectionChanged':false,'rowHotTrackStyle':['dxgvDataRowHover_MaterialCompact',''],'editState':0,'editItemVisibleIndex':-1,'allowSearchFilterTimer':false,'searchPanelFilter':'','allowDelete':false,'allowEdit':false,'allowInsert':false,'columnProp':[[0,,,'nombrePuesto',0,,,,1,,,,,,0],[1,,,'siglasInstitucion',0,,,,3,,,,,,0],[2,,,'vacantes',0,2,,,5,,,,,,0],[3,,,'salario',0,,,,4,,,,,,0],[4,,,'municipio',0,2,,,6,,,,,,0],[5,,,,0,,,,10,,,,,0,0],[6,0,,'nombreInstitucion',0,,,,8,,,,,,0,,1]],'editMode':2,'indentColumnCount':0,'allowChangeColumnHierarchy':false,'allowMultiColumnAutoFilter':false,'adaptiveColumnsOrder':[2,3,1,5,4,0]},null,null,{'adaptiveModeInfo':{'adaptivityMode':2,'hideDataCellsWindowInnerWidth':760,'adaptiveDetailColumnCount':1,'allowTextTruncationInAdaptiveMode':[false,false,false,false,false,false],'adaptiveLayoutColumnIndices':[0,1,3,2,4,5],'allowOnlyOneAdaptiveDetailExpanded':false}});
ASPxClientGridBase.PostponeInitialize('ctl00_MainContent_ultimosEmpleos_gridPuestosPublicados',({'commandButtonIDs':[],'styleInfo':{'sel':{'css':'dxgvSelectedRow_MaterialCompact'},'fi':{'css':'dxgvFocusedRow_MaterialCompact'},'ei':'<tr class="dxgvEditingErrorRow_MaterialCompact">\r\n\t<td class="dxgv" data-colSpan="6" style="border-right-width:0px;"></td>\r\n</tr>','fc':{'css':'dxgvFocusedCell_MaterialCompact'},'bec':{'css':'dxgvBatchEditCell_MaterialCompact dxgv'},'bemc':{'css':'dxgvBatchEditModifiedCell_MaterialCompact dxgv'},'bemergmc':{'css':'dxgvBatchEditModifiedCell_MaterialCompact dxgvBatchEditCell_MaterialCompact dxgv'},'bedi':{'css':'dxgvBatchEditDeletedItem_MaterialCompact dxgv'},'fgi':{'css':'dxgvFocusedGroupRow_MaterialCompact'}}}));

//-->
</script>
                        
            <br />
            &nbsp;&nbsp;<a href="Concursos.aspx">Ver listado completo</a>
            <br />
        </td>
    </tr>
</table>
<br />
            <div class="flex-ayuda">
                <a href="pasos.aspx" target="_self">
                <img alt="¿Cómo participar en un concurso?" src="Content/Images/bannerPasosAbajo.png" id="bannerParticipar" />
                    </a>

                <iframe width="320" height="240" src="https://www.youtube.com/embed/lbAnizGrYvM" frameborder="0" allowfullscreen></iframe>
                
            </div>
        </div>
    </div>


    <div id="footer">
        <div id="footer-wrap">
            <div id="footer-logo"></div>
            <div id="footer-institucion">
            2015 &copy; Copyright Secretaría Técnica y de Planificación de la Presidencia<br />
            <a href="https://www.facebook.com/empleospublicossv/"><i class="fa fa-facebook-square" style="font-size:24px;color:white"></i></a>
            &nbsp;<a href="https://twitter.com/empleopublicosv"><i class="fa fa-twitter-square" style="font-size:24px;color:white"></i></a>
            </div>
            
        </div>
    </div>
</div>
               <div id="ctl00_popupMensaje_PW-1" class="dxpcLite_MaterialCompact dxpclW dxpc-ie" style="z-index:10000;display:none;visibility:hidden;">
	<div class="dxpc-mainDiv dxpc-shadow">
		<div class="dxpc-header" style="padding-left:20px;padding-right:20px;">
			<div class="dxpc-headerContent">
				<span class="dxpc-headerText dx-vam">Mensaje de sistema</span>
			</div><b class="dx-clear"></b>
		</div><div class="dxpc-contentWrapper">
			<div class="dxpc-content" style="padding-left:20px;padding-right:20px;">
				&nbsp;
			</div>
		</div><div class="dxpc-footer">
			
            <div style="width:100%; text-align:center; height:50px;">
                <br />
                     <div class="dxbButton_MaterialCompact edInline dxbButtonSys dxbTSys" id="ctl00_popupMensaje_TPCFm1_btnOk" style="user-select:none;-khtml-user-select:none;-ms-user-select:none;">
				<div class="dxb">
					<input id="ctl00_popupMensaje_TPCFm1_btnOk_I" class="dxb-hb" value="Ok" type="submit" name="ctl00$popupMensaje$TPCFm1$btnOk" /><span class="dx-vam">Ok</span>
				</div>
			</div><script id="dxss_1518735659" type="text/javascript">
<!--
ASPx.AddHoverItems('ctl00_popupMensaje_TPCFm1_btnOk',[[['dxbButtonHover_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddPressedItems('ctl00_popupMensaje_TPCFm1_btnOk',[[['dxbButtonPressed_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddDisabledItems('ctl00_popupMensaje_TPCFm1_btnOk',[[['dxbDisabled_MaterialCompact'],[''],[''],['','TC']]]);
ASPx.AddSelectedItems('ctl00_popupMensaje_TPCFm1_btnOk',[[['dxbf'],[''],['CD']]]);
ASPx.createControl(ASPxClientButton,'ctl00_popupMensaje_TPCFm1_btnOk','btnOk',{'uniqueID':'ctl00$popupMensaje$TPCFm1$btnOk'},{'Click':function(s, e) { popupMensaje.Hide(); } });

//-->
</script>
            </div>
            
		</div>
	</div>
</div><div id="ctl00_popupMensaje_DXPWMB-1" class="dxpcModalBackLite_MaterialCompact" style="z-index:9999;">

</div><table id="ctl00_popupMensaje_LP" class="dxpcLoadingPanel_MaterialCompact dxlpLoadingPanel_MaterialCompact" style="left:0px;top:0px;z-index:30000;display:none;">
	<tr>
		<td class="dx" style="padding-right:0px;"><img class="dxlp-loadingImage dxlp-imgPosLeft" src="/DXR.axd?r=1_58-MVpNf" alt="" style="vertical-align:middle;" /></td><td class="dx" style="padding-left:0px;"><span id="ctl00_popupMensaje_TL">Cargando&hellip;</span></td>
	</tr>
</table><div id="ctl00_popupMensaje_LD" class="dxpcLoadingDiv_MaterialCompact dxlpLoadingDiv_MaterialCompact dx-ft" style="left:0px;top:0px;z-index:29999;display:none;position:absolute;">

</div><script id="dxss_1562554604" type="text/javascript">
<!--
ASPx.createControl(ASPxClientPopupControl,'ctl00_popupMensaje','popupMensaje',{'encodeHtml':false,'callBack':function(arg) { WebForm_DoCallback('ctl00$popupMensaje',arg,ASPx.Callback,'ctl00_popupMensaje',ASPx.CallbackError,true); },'uniqueID':'ctl00$popupMensaje','popupAnimationType':'fade','closeAnimationType':'fade','popupHorizontalAlign':'WindowCenter','popupVerticalAlign':'WindowCenter','isPopupPositionCorrectionOn':false,'modal':true,'width':400,'widthFromServer':true,'SSLSecureBlankUrl':'/DXR.axd?r=1_0-MVpNf'});

//-->
</script>
    </form>
</body>
</html>