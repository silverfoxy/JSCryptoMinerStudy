<!doctype html><html lang="es"><head prefix="og: http://ogp.me/ns#"><meta charset="UTF-8"><title>Radios de El Salvador en linea, emisoras de El Salvador online</title><meta name="description" content="Todas las radios El Salvador en sólo una página. Súper fácil y 100% gratis."><meta name="theme-color" content="#002029"><meta name="viewport" content="width=device-width, initial-scale=1.0"><meta property="fb:admins" content="100002936790534"><meta property="og:locale" content="es_LA"><meta property="og:url" content="http://www.radios.com.sv/"><meta property="og:title" content="Radios de El Salvador en linea, emisoras de El Salvador online"><meta property="og:site_name" content="Radios.com.sv"><meta property="og:description" content="Todas las radios El Salvador en sólo una página. Súper fácil y 100% gratis."><meta property="og:image" content="https://cdn.webrad.io/images/countries/el-salvador-logo_512x512.png"><meta property="og:type" content="website"><link rel="canonical" href="http://www.radios.com.sv/"><link rel="dns-prefetch" href="//api.webrad.io"><link rel="dns-prefetch" href="//apis.google.com"><link rel="dns-prefetch" href="//cdn.trackjs.com"><link rel="dns-prefetch" href="//cdn.webrad.io"><link rel="dns-prefetch" href="//cdnjs.cloudflare.com"><link rel="dns-prefetch" href="//connect.facebook.net"><link rel="dns-prefetch" href="//pagead2.googlesyndication.com"><link rel="dns-prefetch" href="//platform.twitter.com"><link rel="dns-prefetch" href="//webrad.io"><link rel="dns-prefetch" href="//www.googletagmanager.com"><link rel="preconnect" href="//api.webrad.io"><link rel="preconnect" href="//apis.google.com"><link rel="preconnect" href="//cdn.trackjs.com"><link rel="preconnect" href="//cdn.webrad.io"><link rel="preconnect" href="//cdnjs.cloudflare.com"><link rel="preconnect" href="//connect.facebook.net"><link rel="preconnect" href="//pagead2.googlesyndication.com"><link rel="preconnect" href="//platform.twitter.com"><link rel="preconnect" href="//www.googletagmanager.com"><link rel="prefetch" href="https://cdn.webrad.io/images/icon-error.png"><link rel="prefetch" href="https://cdn.webrad.io/images/icon-flash.png"><link rel="prefetch" href="https://cdn.webrad.io/images/icon-open.png"><link rel="prefetch" href="https://cdn.webrad.io/images/icon-play.png"><link rel="prefetch" href="https://cdn.webrad.io/images/icon-sound-off.png"><link rel="prefetch" href="https://cdnjs.cloudflare.com/ajax/libs/cookieconsent2/3.0.6/cookieconsent.min.css"><link rel="prefetch" href="https://cdnjs.cloudflare.com/ajax/libs/cookieconsent2/3.0.6/cookieconsent.min.js"><link rel="prefetch" href="https://cdnjs.cloudflare.com/ajax/libs/dashjs/2.6.6/dash.mediaplayer.min.js"><link rel="prefetch" href="https://cdnjs.cloudflare.com/ajax/libs/hls.js/0.8.9/hls.light.min.js"><link rel="preload" href="https://cdn.webrad.io/images/icon-load.gif" as="image"><link rel="preload" href="https://cdn.webrad.io/images/icon-sound-on.png" as="image"><link rel="preload" href="https://cdn.webrad.io/images/icon-stop.png" as="image"><link rel="preload" href="http://api.webrad.io/data/streams/36/scan-96-1-fm" as="fetch" type="application/json" crossorigin><link rel="preload" href="https://cdn.webrad.io/fonts/icomoon.ttf" as="font" type="font/ttf" crossorigin="anonymous"><link rel="preload" href="https://cdn.webrad.io/js/jquery.main-4.0.16.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdn.webrad.io/js/jquery.mobilenav.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdn.webrad.io/js/jquery.openclose.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/algoliasearch/3.24.12/algoliasearchLite.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/bowser/1.9.2/bowser.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/hogan.js/3.0.2/hogan.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/jquery/3.3.1/jquery.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/rangeslider.js/2.3.2/rangeslider.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/simplebar/2.5.1/simplebar.min.js" as="script" crossorigin="anonymous"><link rel="preload" href="https://cdnjs.cloudflare.com/ajax/libs/soundmanager2/2.97a.20170601/script/soundmanager2-nodebug-jsmin.js" as="script" crossorigin="anonymous"><link rel="shortcut icon" href="https://cdn.webrad.io/images/countries/el-salvador.ico"><link rel="stylesheet" href="https://cdn.webrad.io/css/main-4.0.6.min.css"><script>window._trackJs={console:{display:!1},enabled:8E-4>Math.random()?!0:!1,token:"73faad723c2e459eafb494db926fccb4",version:"4.0.16"};window.SM2_DEFER=!0;var webradioConfig={countryCode:"SV",debugMode:0,domainID:36,languageCode:"es",slugDomain:"radios-com-sv",urlApi:"http://api.webrad.io/",urlStatic:"https://cdn.webrad.io/",cookieConsent:{version:"3.0.6",link:"Info",href:"/politica-de-privacidad/"},algolia:[{"applicationId":"3ZTZWUB3YF","apiKey":"69c38d1d7696f10303d883840d265170"}],dashJs:{version:"2.6.6"},facebook:{countryCode:"LA",version:"2.12"},hlsJs:{version:"0.8.9"},txt:{cookie:"Este sitio web utiliza cookies para asegurarse de que puedas aprovechar al m\u00e1ximo tu experiencia en nuestro sitio web",error:"Error",loading:"Cargando",mute:"Desactivar o reactivar audio",no_audio:"Sin audio durante m\u00e1s de un mes, lo comprobamos semanalmente",ok:"OK",play:"Sonar",popup:"Escuchar aqui",search_for:"Resultados de la b\u00fasqueda de %s",search_none:"No hay resultados para %s",start:"Inicio",stop:"Parar",volume:"Control de volumen"}};</script><script src="https://pagead2.googlesyndication.com/pagead/js/adsbygoogle.js" async></script><script src="https://www.googletagmanager.com/gtag/js?id=UA-43921502-1" async></script><script src="https://cdn.trackjs.com/releases/current/tracker.js" async crossorigin="anonymous"></script><script>window.dataLayer=window.dataLayer||[];function gtag(){dataLayer.push(arguments)}gtag("js",new Date);gtag("config","UA-43921502-1",{cookie_domain:"radios.com.sv"});setTimeout(function(){gtag("event","60 seconds",{event_category:"Read"})},6E4);</script></head><body class="ltr"><div id="wrapper">
	<header id="header">
		<div class="top-header"><div class="container"><a class="country-opener" href="http://www.radios.com.sv/" title="El Salvador"><img src="https://cdn.webrad.io/images/countries/el-salvador_14x11.png" alt="El Salvador" height="11" width="14"></a><div class="nav-holder"><ul class="country-list"><li><a href="http://www.radioarg.com/" title="Argentina"><img src="https://cdn.webrad.io/images/countries/argentina_14x11.png" alt="Argentina" height="11" width="14"></a></li><li><a href="http://www.radios.com.bo/" title="Bolivia"><img src="https://cdn.webrad.io/images/countries/bolivia_14x11.png" alt="Bolivia" height="11" width="14"></a></li><li><a href="http://www.radiosaovivo.net/" title="Brasil"><img src="https://cdn.webrad.io/images/countries/brazil_14x11.png" alt="Brasil" height="11" width="14"></a></li><li><a href="http://www.emisora.cl/" title="Chile"><img src="https://cdn.webrad.io/images/countries/chile_14x11.png" alt="Chile" height="11" width="14"></a></li><li><a href="http://www.radios.com.co/" title="Colombia"><img src="https://cdn.webrad.io/images/countries/colombia_14x11.png" alt="Colombia" height="11" width="14"></a></li><li><a href="http://www.radios.co.cr/" title="Costa Rica"><img src="https://cdn.webrad.io/images/countries/costa-rica_14x11.png" alt="Costa Rica" height="11" width="14"></a></li><li><a href="http://www.radiosdecuba.com/" title="Cuba"><img src="https://cdn.webrad.io/images/countries/cuba_14x11.png" alt="Cuba" height="11" width="14"></a></li><li><a href="http://www.radios.com.do/" title="República Dominicana"><img src="https://cdn.webrad.io/images/countries/dominican-republic_14x11.png" alt="República Dominicana" height="11" width="14"></a></li><li><a href="http://www.radios.com.ec/" title="Ecuador"><img src="https://cdn.webrad.io/images/countries/ecuador_14x11.png" alt="Ecuador" height="11" width="14"></a></li><li><a href="http://www.emisoras.com.gt/" title="Guatemala"><img src="https://cdn.webrad.io/images/countries/guatemala_14x11.png" alt="Guatemala" height="11" width="14"></a></li><li><a href="http://www.radio.ht/" title="Haïti"><img src="https://cdn.webrad.io/images/countries/haiti_14x11.png" alt="Haïti" height="11" width="14"></a></li><li><a href="http://www.radios.hn/" title="Honduras"><img src="https://cdn.webrad.io/images/countries/honduras_14x11.png" alt="Honduras" height="11" width="14"></a></li><li><a href="http://www.jamaicaradio.net/" title="Jamaica"><img src="https://cdn.webrad.io/images/countries/jamaica_14x11.png" alt="Jamaica" height="11" width="14"></a></li><li><a href="http://www.emisoras.com.mx/" title="México"><img src="https://cdn.webrad.io/images/countries/mexico_14x11.png" alt="México" height="11" width="14"></a></li><li><a href="http://www.radios.co.ni/" title="Nicaragua"><img src="https://cdn.webrad.io/images/countries/nicaragua_14x11.png" alt="Nicaragua" height="11" width="14"></a></li><li><a href="http://www.radios.com.pa/" title="Panamá"><img src="https://cdn.webrad.io/images/countries/panama_14x11.png" alt="Panamá" height="11" width="14"></a></li><li><a href="http://www.emisoras.com.py/" title="Paraguay"><img src="https://cdn.webrad.io/images/countries/paraguay_14x11.png" alt="Paraguay" height="11" width="14"></a></li><li><a href="http://www.radios.com.pe/" title="Perú"><img src="https://cdn.webrad.io/images/countries/peru_14x11.png" alt="Perú" height="11" width="14"></a></li><li><a href="http://www.radiosdepuertorico.com/" title="Puerto Rico"><img src="https://cdn.webrad.io/images/countries/puerto-rico_14x11.png" alt="Puerto Rico" height="11" width="14"></a></li><li><a href="http://www.surinaamseradio.com/" title="Suriname"><img src="https://cdn.webrad.io/images/countries/suriname_14x11.png" alt="Suriname" height="11" width="14"></a></li><li><a href="http://www.trinidadradiostations.net/" title="Trinidad and Tobago"><img src="https://cdn.webrad.io/images/countries/trinidad-and-tobago_14x11.png" alt="Trinidad and Tobago" height="11" width="14"></a></li><li><a href="http://www.radios.com.uy/" title="Uruguay"><img src="https://cdn.webrad.io/images/countries/uruguay_14x11.png" alt="Uruguay" height="11" width="14"></a></li><li><a href="http://www.radios.co.ve/" title="Venezuela"><img src="https://cdn.webrad.io/images/countries/venezuela_14x11.png" alt="Venezuela" height="11" width="14"></a></li></ul><a class="more" href="http://www.radiowebsites.org/" title="Más países">Más países</a></div></div></div>		<div class="container">
			<div class="logo"><a href="http://www.radios.com.sv/"><img class="ico" src="https://cdn.webrad.io/images/equalizer.gif" alt="Radios.com.sv" height="14" width="23">Radios<span>.com.sv</span></a></div><div class="add-box-top"><ins class="adsbygoogle" data-ad-client="ca-pub-6771940464972938" data-ad-slot="4118848263" data-ad-format="auto"></ins><script>(adsbygoogle=window.adsbygoogle||[]).push({});</script></div>		</div>
	</header>
	<main id="main">
		<div class="container">
			<section id="content">
				<div class="content-holder">
					<div class="head"><a class="menu-opener" href="#"><span>Menú</span></a><form class="search-form" action="#"><div class="input-holder"><button type="submit" aria-label="Buscar" name="Buscar"><i class="icon-search"></i></button><input type="search" id="search-input-head" aria-label="Buscar" autocomplete="on" placeholder="Buscar" required spellcheck="false"></div></form><div class="social-links"><div id="fb-root"></div><div class="social-btn fb-like" data-href="http://www.radios.com.sv/" data-layout="button_count" data-width="150"></div><div class="social-btn"><div class="g-plusone" data-href="http://www.radios.com.sv/" data-size="medium"></div></div><a class="social-btn twitter-share-button" href="https://twitter.com/share?url=http%3A%2F%2Fwww.radios.com.sv%2F&amp;via=emisoraselsalva&amp;text=Estoy+disfrutando+de+las+estaciones+de+radio+de+El+Salvador+en&amp;count=horizontal&amp;lang=es" title="Twitter"></a></div></div><span class="overlay"></span><div class="menu-area" data-simplebar><form class="search-form" action="#"><div class="input-holder"><button type="submit" aria-label="Buscar" name="Buscar"><i class="icon-search"></i></button><input type="search" id="search-input-menu" aria-label="Buscar" autocomplete="on" placeholder="Buscar cualquier emisora de radio" required spellcheck="false"></div></form><div class="box active"><strong class="title"><a class="opener" href="#">Géneros</a></strong><a class="more" href="http://www.radios.com.sv/generos/">Todos los géneros</a><div class="slide"><ul class="menu-list"><li><a href="http://www.radios.com.sv/genero/musica-mundial/">Música Mundial</a></li><li><a href="http://www.radios.com.sv/genero/top-40/">Top 40</a></li><li><a href="http://www.radios.com.sv/genero/religion/">Religión</a></li><li><a href="http://www.radios.com.sv/genero/musica-latina/">Música Latina</a></li><li><a href="http://www.radios.com.sv/genero/cristiano/">Cristiano</a></li><li><a href="http://www.radios.com.sv/genero/entrevistas/">Entrevistas</a></li><li><a href="http://www.radios.com.sv/genero/espiritualidad/">Espiritualidad</a></li><li><a href="http://www.radios.com.sv/genero/noticias/">Noticias</a></li><li><a href="http://www.radios.com.sv/genero/contemporaneo/">Contemporáneo</a></li><li><a href="http://www.radios.com.sv/genero/crist-espanol/">Crist. Español</a></li></ul></div></div><div class="box active"><strong class="title"><a class="opener" href="#">Regiones</a></strong><div class="slide"><ul class="menu-list"><li><a href="http://www.radios.com.sv/region/san-salvador-1/">San Salvador 1</a></li><li><a href="http://www.radios.com.sv/region/san-salvador-2/">San Salvador 2</a></li><li><a href="http://www.radios.com.sv/region/otras-regiones-1/">Otras regiones 1</a></li><li><a href="http://www.radios.com.sv/region/otras-regiones-2/">Otras regiones 2</a></li></ul></div></div><div class="box active"><strong class="title"><a class="opener" href="#">Frecuencias</a></strong><div class="slide"><ul class="menu-list"><li><a href="http://www.radios.com.sv/bautista/" title="Radio Bautista 89.7 FM">89.7 FM</a></li><li><a href="http://www.radios.com.sv/la-caliente/" title="La Caliente San Miguel 90.1 FM">90.1 FM</a></li><li><a href="http://www.radios.com.sv/exa/" title="Exa 91.3 FM">91.3 FM</a></li><li><a href="http://www.radios.com.sv/doremix/" title="Radio Doremix 92.5 FM">92.5-1 FM</a></li><li><a href="http://www.radios.com.sv/club/" title="Radio Club 92.5 FM">92.5-2 FM</a></li><li><a href="http://www.radios.com.sv/laser/" title="Radio Laser 92.9 FM">92.9 FM</a></li><li><a href="http://www.radios.com.sv/globo/" title="FM Globo 93.3">93.3 FM</a></li><li><a href="http://www.radios.com.sv/el-mundo/" title="Radio el Mundo 93.7 FM">93.7 FM</a></li><li><a href="http://www.radios.com.sv/fabulosa-santa-rosa-de-lima/" title="Radio La Fabulosa 94.1 FM Santa Rosa de Lima">94.1 FM</a></li><li><a href="http://www.radios.com.sv/vox/" title="Vox 94.5 FM">94.5 FM</a></li><li><a href="http://www.radios.com.sv/coco/" title="Radio Coco 94.9 FM">94.9-1 FM</a></li><li><a href="http://www.radios.com.sv/astral/" title="Radio Astral 94.9 FM">94.9-2 FM</a></li><li><a href="http://www.radios.com.sv/galaxia/" title="Radio Galaxia 94.9 FM">94.9-3 FM</a></li><li><a href="http://www.radios.com.sv/eco/" title="Radio Eco 95.3 FM">95.3-1 FM</a></li><li><a href="http://www.radios.com.sv/kyrios/" title="Radio Kyrios 95.3 FM">95.3-2 FM</a></li><li><a href="http://www.radios.com.sv/verdad/" title="Radio Verdad 95.7 FM">95.7 FM</a></li><li><a href="http://www.radios.com.sv/scan/" title="Scan 96.1 FM">96.1 FM</a></li><li><a href="http://www.radios.com.sv/adventista/" title="Radio Adventista 96.5 FM">96.5-1 FM</a></li><li><a href="http://www.radios.com.sv/agape/" title="Agape Radio Oriente 96.5 FM">96.5-2 FM</a></li><li><a href="http://www.radios.com.sv/nacional/" title="Radio Nacional El Salvador">96.9 FM</a></li><li><a href="http://www.radios.com.sv/luz/" title="Radio Luz 97.7 FM">97.7 FM</a></li><li><a href="http://www.radios.com.sv/pantera-san-salvador/" title="Radio La Pantera 98.1 FM San Salvador">98.1 FM</a></li><li><a href="http://www.radios.com.sv/cadena-cuscatlan/" title="Radio Cadena Cuscatlán">98.5 FM</a></li><li><a href="http://www.radios.com.sv/la-mejor/" title="La Mejor 98.9 FM">98.9 FM</a></li><li><a href="http://www.radios.com.sv/mesias/" title="Radio Mesías 99.3 FM">99.3 FM</a></li><li><a href="http://www.radios.com.sv/rx/" title="Radio RX FM 99.7">99.7-1 FM</a></li><li><a href="http://www.radios.com.sv/full/" title="Radio Full online 99.7 FM">99.7-2 FM</a></li><li><a href="http://www.radios.com.sv/abc/" title="ABC 100.1 FM Stereo">100.1 FM</a></li><li><a href="http://www.radios.com.sv/radio-la-chevere/" title="Radio La Chévere 100.9 FM">100.9 FM</a></li><li><a href="http://www.radios.com.sv/monumental/" title="Radio Monumental 101.3 FM">101.3 FM</a></li><li><a href="http://www.radios.com.sv/femenina/" title="Femenina 102.5 FM">102.5 FM</a></li><li><a href="http://www.radios.com.sv/nueve/" title="Radio 102.9 FM">102.9 FM</a></li><li><a href="http://www.radios.com.sv/clasica/" title="Clásica Online 103.3 FM">103.3 FM</a></li><li><a href="http://www.radios.com.sv/yskl/" title="Radio YSKL 104.1 FM">104.1 FM</a></li><li><a href="http://www.radios.com.sv/radio-fiesta/" title="Radio Fiesta 104.9 FM">104.9 FM</a></li><li><a href="http://www.radios.com.sv/soda-stereo/" title="Soda Stereo 105.3 FM">105.3 FM</a></li><li><a href="http://www.radios.com.sv/yxy/" title="Radio YXY 105.7 FM">105.7 FM</a></li><li><a href="http://www.radios.com.sv/el-camino/" title="El Camino 106.1 FM">106.1-1 FM</a></li><li><a href="http://www.radios.com.sv/impacto/" title="Radio Impacto 106.1 FM">106.1-2 FM</a></li><li><a href="http://www.radios.com.sv/ranchera/" title="Ranchera 106.5 FM">106.5 FM</a></li><li><a href="http://www.radios.com.sv/mi-gente/" title="Radio Cadena Mi Gente">700 AM</a></li><li><a href="http://www.radios.com.sv/chaparrastique/" title="Radio Chaparrastique 106.1 FM">950 AM</a></li><li><a href="http://www.radios.com.sv/getsemani-la-union/" title="Radio Getsemani 1390 AM La Unión">1390 AM</a></li></ul></div></div></div><div id="search-results"></div>					<div class="radio-section" id="content-area">
						<h2>Radios de El Salvador</h2>
						<div id="radio"><div class="loading" id="radio-track"><div class="left-box"><div class="img-box"><img id="radio-logo" src="https://cdn.webrad.io/images/spacer.gif" alt="" height="66" width="96"></div><div class="text-box"><strong class="title" id="radio-title"></strong><span class="fm-text" id="radio-frequency"></span></div></div><div class="btn-holder"><a class="btn white" id="radio-link" href="#" rel="nofollow noopener" target="_blank">Web</a><a class="btn white" id="radio-no-audio" href="http://www.radios.com.sv/ayuda/" rel="nofollow noopener" target="_blank">¿No funciona?</a></div></div><div class="radio-player"><div class="loading" id="radio-controls"><span class="btn-play"></span><span class="ico-load"></span><span class="rangeslider"></span></div></div></div><ul id="radios"><li class="item-1"><span><a href="http://www.radios.com.sv/#scan-96-1-fm" title="Scan 96.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/scan-96-1-fm.png" alt="Scan 96.1 FM" height="66" width="96"></a></span></li><li class="item-2"><span><a href="http://www.radios.com.sv/#radio-la-chevere-100-9-fm" title="Radio La Chévere 100.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-la-chevere-100-9-fm.png" alt="Radio La Chévere 100.9 FM" height="66" width="96"></a></span></li><li class="item-3"><span><a href="http://www.radios.com.sv/#radio-fiesta-104-9-fm" title="Radio Fiesta 104.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-fiesta-104-9-fm.png" alt="Radio Fiesta 104.9 FM" height="66" width="96"></a></span></li><li class="item-4"><span><a href="http://www.radios.com.sv/#ranchera-106-5-fm" title="Ranchera 106.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/ranchera-106-5-fm.png" alt="Ranchera 106.5 FM" height="66" width="96"></a></span></li><li class="item-5"><span><a href="http://www.radios.com.sv/#radio-yskl-104-1-fm" title="Radio YSKL 104.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-yskl-104-1-fm.png" alt="Radio YSKL 104.1 FM" height="66" width="96"></a></span></li><li class="item-6"><span><a href="http://www.radios.com.sv/#radio-getsemani-1390-am-la-union" title="Radio Getsemani 1390 AM La Unión"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-getsemani-1390-am-la-union.png" alt="Radio Getsemani 1390 AM La Unión" height="66" width="96"></a></span></li><li class="item-7"><span><a href="http://www.radios.com.sv/#radio-monumental-101-3-fm" title="Radio Monumental 101.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-monumental-101-3-fm.png" alt="Radio Monumental 101.3 FM" height="66" width="96"></a></span></li><li class="item-8"><span><a href="http://www.radios.com.sv/#radio-yxy-105-7-fm" title="Radio YXY 105.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-yxy-105-7-fm.png" alt="Radio YXY 105.7 FM" height="66" width="96"></a></span></li><li class="item-9"><span><a href="http://www.radios.com.sv/#la-mejor-98-9-fm" title="La Mejor 98.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/la-mejor-98-9-fm.png" alt="La Mejor 98.9 FM" height="66" width="96"></a></span></li><li class="item-10"><span><a href="http://www.radios.com.sv/#fm-globo-93-3" title="FM Globo 93.3"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/fm-globo-93-3.png" alt="FM Globo 93.3" height="66" width="96"></a></span></li><li class="item-11"><span><a href="http://www.radios.com.sv/#radio-la-pantera-98-1-fm-san-salvador" title="Radio La Pantera 98.1 FM San Salvador"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-la-pantera-98-1-fm-san-salvador.png" alt="Radio La Pantera 98.1 FM San Salvador" height="66" width="96"></a></span></li><li class="item-12"><span><a href="http://www.radios.com.sv/#radio-cadena-cuscatlan" title="Radio Cadena Cuscatlán"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-cadena-cuscatlan.png" alt="Radio Cadena Cuscatlán" height="66" width="96"></a></span></li><li class="item-13"><span><a href="http://www.radios.com.sv/#vox-94-5-fm" title="Vox 94.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/vox-94-5-fm.png" alt="Vox 94.5 FM" height="66" width="96"></a></span></li><li class="item-14"><span><a href="http://www.radios.com.sv/#radio-cadena-mi-gente" title="Radio Cadena Mi Gente"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-cadena-mi-gente.png" alt="Radio Cadena Mi Gente" height="66" width="96"></a></span></li><li class="item-15"><span><a href="http://www.radios.com.sv/#femenina-102-5-fm" title="Femenina 102.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/femenina-102-5-fm.png" alt="Femenina 102.5 FM" height="66" width="96"></a></span></li><li class="item-16"><span><a href="http://www.radios.com.sv/#radio-eco-95-3-fm" title="Radio Eco 95.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-eco-95-3-fm.png" alt="Radio Eco 95.3 FM" height="66" width="96"></a></span></li><li class="item-17"><span><a href="http://www.radios.com.sv/#exa-91-3-fm" title="Exa 91.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/exa-91-3-fm.png" alt="Exa 91.3 FM" height="66" width="96"></a></span></li><li class="item-18"><span><a href="http://www.radios.com.sv/#radio-club-92-5-fm" title="Radio Club 92.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-club-92-5-fm.png" alt="Radio Club 92.5 FM" height="66" width="96"></a></span></li><li class="item-19"><span><a href="http://www.radios.com.sv/#radio-impacto-106-1-fm" title="Radio Impacto 106.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-impacto-106-1-fm.png" alt="Radio Impacto 106.1 FM" height="66" width="96"></a></span></li><li class="item-20"><span><a href="http://www.radios.com.sv/#radio-chaparrastique-106-1-fm" title="Radio Chaparrastique 106.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-chaparrastique-106-1-fm.png" alt="Radio Chaparrastique 106.1 FM" height="66" width="96"></a></span></li><li class="item-21"><span><a href="http://www.radios.com.sv/#radio-luz-97-7-fm" title="Radio Luz 97.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-luz-97-7-fm.png" alt="Radio Luz 97.7 FM" height="66" width="96"></a></span></li><li class="item-22"><span><a href="http://www.radios.com.sv/#radio-coco-94-9-fm" title="Radio Coco 94.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-coco-94-9-fm.png" alt="Radio Coco 94.9 FM" height="66" width="96"></a></span></li><li class="item-23"><span><a href="http://www.radios.com.sv/#radio-doremix-92-5-fm" title="Radio Doremix 92.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-doremix-92-5-fm.png" alt="Radio Doremix 92.5 FM" height="66" width="96"></a></span></li><li class="item-24"><span><a href="http://www.radios.com.sv/#radio-rx-fm-99-7" title="Radio RX FM 99.7"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-rx-fm-99-7.png" alt="Radio RX FM 99.7" height="66" width="96"></a></span></li><li class="item-25"><span><a href="http://www.radios.com.sv/#clasica-online-103-3-fm" title="Clásica Online 103.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/clasica-online-103-3-fm.png" alt="Clásica Online 103.3 FM" height="66" width="96"></a></span></li><li class="item-26"><span><a href="http://www.radios.com.sv/#radio-bautista-89-7-fm" title="Radio Bautista 89.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-bautista-89-7-fm.png" alt="Radio Bautista 89.7 FM" height="66" width="96"></a></span></li><li class="item-27"><span><a href="http://www.radios.com.sv/#radio-astral-94-9-fm" title="Radio Astral 94.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-astral-94-9-fm.png" alt="Radio Astral 94.9 FM" height="66" width="96"></a></span></li><li class="item-28"><span><a href="http://www.radios.com.sv/#radio-102-9-fm" title="Radio 102.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-102-9-fm.png" alt="Radio 102.9 FM" height="66" width="96"></a></span></li><li class="item-29"><span><a href="http://www.radios.com.sv/#radio-mesias-99-3-fm" title="Radio Mesías 99.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-mesias-99-3-fm.png" alt="Radio Mesías 99.3 FM" height="66" width="96"></a></span></li><li class="item-30"><span><a href="http://www.radios.com.sv/#radio-full-online-99-7-fm" title="Radio Full online 99.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-full-online-99-7-fm.png" alt="Radio Full online 99.7 FM" height="66" width="96"></a></span></li><li class="item-31"><span><a href="http://www.radios.com.sv/#abc-100-1-fm-stereo" title="ABC 100.1 FM Stereo"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/abc-100-1-fm-stereo.png" alt="ABC 100.1 FM Stereo" height="66" width="96"></a></span></li><li class="item-32"><span><a href="http://www.radios.com.sv/#radio-el-mundo-93-7-fm" title="Radio el Mundo 93.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-el-mundo-93-7-fm.png" alt="Radio el Mundo 93.7 FM" height="66" width="96"></a></span></li><li class="item-33"><span><a href="http://www.radios.com.sv/#radio-verdad-95-7-fm" title="Radio Verdad 95.7 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-verdad-95-7-fm.png" alt="Radio Verdad 95.7 FM" height="66" width="96"></a></span></li><li class="item-34"><span><a href="http://www.radios.com.sv/#el-camino-106-1-fm" title="El Camino 106.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/el-camino-106-1-fm.png" alt="El Camino 106.1 FM" height="66" width="96"></a></span></li><li class="item-35"><span><a href="http://www.radios.com.sv/#radio-laser-92-9-fm" title="Radio Laser 92.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-laser-92-9-fm.png" alt="Radio Laser 92.9 FM" height="66" width="96"></a></span></li><li class="item-36"><span><a href="http://www.radios.com.sv/#radio-galaxia-94-9-fm" title="Radio Galaxia 94.9 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-galaxia-94-9-fm.png" alt="Radio Galaxia 94.9 FM" height="66" width="96"></a></span></li><li class="item-37"><span><a href="http://www.radios.com.sv/#radio-adventista-96-5-fm" title="Radio Adventista 96.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-adventista-96-5-fm.png" alt="Radio Adventista 96.5 FM" height="66" width="96"></a></span></li><li class="item-38"><span><a href="http://www.radios.com.sv/#radio-kyrios-95-3-fm" title="Radio Kyrios 95.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-kyrios-95-3-fm.png" alt="Radio Kyrios 95.3 FM" height="66" width="96"></a></span></li><li class="item-39"><span><a href="http://www.radios.com.sv/#agape-radio-oriente-96-5-fm" title="Agape Radio Oriente 96.5 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/agape-radio-oriente-96-5-fm.png" alt="Agape Radio Oriente 96.5 FM" height="66" width="96"></a></span></li><li class="item-40"><span><a href="http://www.radios.com.sv/#la-caliente-san-miguel-90-1-fm" title="La Caliente San Miguel 90.1 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/la-caliente-san-miguel-90-1-fm.png" alt="La Caliente San Miguel 90.1 FM" height="66" width="96"></a></span></li><li class="item-41"><span><a href="http://www.radios.com.sv/#radio-la-fabulosa-94-1-fm-santa-rosa-de-lima" title="Radio La Fabulosa 94.1 FM Santa Rosa de Lima"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-la-fabulosa-94-1-fm-santa-rosa-de-lima.png" alt="Radio La Fabulosa 94.1 FM Santa Rosa de Lima" height="66" width="96"></a></span></li><li class="item-42"><span><a href="http://www.radios.com.sv/#soda-stereo-105-3-fm" title="Soda Stereo 105.3 FM"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/soda-stereo-105-3-fm.png" alt="Soda Stereo 105.3 FM" height="66" width="96"></a></span></li><li class="item-43"><span><a href="http://www.radios.com.sv/#radio-nacional-el-salvador" title="Radio Nacional El Salvador"><img class="cover" src="https://cdn.webrad.io/images/logos/radios-com-sv/radio-nacional-el-salvador.png" alt="Radio Nacional El Salvador" height="66" width="96"></a></span></li></ul>					</div>
				</div>
				<div class="add-box-bottom"><ins class="adsbygoogle" data-ad-client="ca-pub-6771940464972938" data-ad-slot="9819511909" data-ad-format="auto"></ins><script>(adsbygoogle=window.adsbygoogle||[]).push({});</script></div>			</section>
			<div class="add-box-side"><ins class="adsbygoogle" data-ad-client="ca-pub-6771940464972938" data-ad-slot="4310419956" data-ad-format="auto"></ins><script>(adsbygoogle=window.adsbygoogle||[]).push({});</script></div>		</div>
	</main>
	<footer id="footer">
		<div class="container">
			<ul class="socialnetworks"><li><a class="icon-facebook" href="https://www.facebook.com/Emisoras.de.El.Salvador/" rel="nofollow noopener" target="_blank" title="Facebook"></a></li><li><a class="icon-google-plus" href="https://plus.google.com/104320019291459551754" rel="nofollow noopener" target="_blank" title="Google+"></a></li><li><a class="icon-twitter" href="https://twitter.com/emisoraselsalva" rel="nofollow noopener" target="_blank" title="Twitter"></a></li></ul><ul class="footer-nav"><li><a href="http://www.radios.com.sv/incluir-tu-radio/" rel="nofollow">Incluir tu radio</a></li><li><a href="http://www.radios.com.sv/ayuda/" rel="nofollow">Ayuda</a></li><li><a href="http://www.radios.com.sv/region/nuevo/" rel="nofollow">Nuevo</a></li><li><a href="http://www.radios.com.sv/politica-de-privacidad/" rel="nofollow">Política de privacidad</a></li><li><a href="mailto:info@radios.com.sv">Contáctenos</a></li><li><a href="http://www.radios.com.sv/dmca/" rel="nofollow">DMCA</a></li></ul>		</div>
	</footer>
</div>
<script src="https://cdnjs.cloudflare.com/ajax/libs/algoliasearch/3.24.12/algoliasearchLite.min.js" crossorigin="anonymous"></script><script src="https://cdnjs.cloudflare.com/ajax/libs/bowser/1.9.2/bowser.min.js" crossorigin="anonymous"></script><script src="https://cdnjs.cloudflare.com/ajax/libs/hogan.js/3.0.2/hogan.min.js" crossorigin="anonymous"></script><script src="https://cdnjs.cloudflare.com/ajax/libs/jquery/3.3.1/jquery.min.js" crossorigin="anonymous"></script><script src="https://cdn.webrad.io/js/jquery.mobilenav.min.js" crossorigin="anonymous"></script><script src="https://cdn.webrad.io/js/jquery.openclose.min.js" crossorigin="anonymous"></script><script src="https://cdnjs.cloudflare.com/ajax/libs/rangeslider.js/2.3.2/rangeslider.min.js" crossorigin="anonymous"></script><script src="https://cdnjs.cloudflare.com/ajax/libs/soundmanager2/2.97a.20170601/script/soundmanager2-nodebug-jsmin.js" crossorigin="anonymous"></script><script src="https://cdn.webrad.io/js/jquery.main-4.0.16.min.js" crossorigin="anonymous"></script><!--[if lte IE 9]><script src="https://cdnjs.cloudflare.com/ajax/libs/jquery-ajaxtransport-xdomainrequest/1.0.4/jquery.xdomainrequest.min.js" crossorigin="anonymous"></script><![endif]--><!--[if (gt IE 9)|!(IE)]><!--><script src="https://cdnjs.cloudflare.com/ajax/libs/simplebar/2.5.1/simplebar.min.js" async crossorigin="anonymous"></script><!--<![endif]--></body></html>