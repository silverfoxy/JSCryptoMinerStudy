<!DOCTYPE html>
<!-- Open Html -->
<html lang="es-ES" prefix="og: http://ogp.me/ns#">
	<!-- Open Head -->
	<head>

<div class="container" >
<div class="row " style="margin-left: -5px; z-index:1000; position:absolute width:100px;">
		<div class="col-md-12 col-lg-12 hidden-xs hidden-sm " style="color: #FFF; width:100px; margin-top: 1px; z-index:1000; position:absolute">
<img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/UNICAES_New_Logo_08.jpg" width="67"></img>

</div>
</div>
</div>
		<meta charset="UTF-8"/>

<meta name="viewport" content="width=device-width, initial-scale=1, maximum-scale=1">
<meta name="google-site-verification" content="o6je6KcS68eAXTCx8vREM6I3ULzxSEQ4l5bnHnUNHBk" />






<!--[if lt IE 9]>
<script src="https://oss.maxcdn.com/html5shiv/3.7.2/html5shiv.min.js"></script>
<script src="https://oss.maxcdn.com/respond/1.4.2/respond.min.js"></script>
<script src="http://css3-mediaqueries-js.googlecode.com/svn/trunk/css3-mediaqueries.js"></script>
<![endif]--><title>Universidad Católica de El Salvador - UNICAES</title>

<!-- This site is optimized with the Yoast SEO Premium plugin v6.2 - https://yoa.st/1yg?utm_content=6.2 -->
<meta name="description" content="La UNICAES es una Institución de educación superior que forma profesionales integrales, con principios cristianos y conocimientos técnicos y científicos"/>
<link rel="canonical" href="http://www.catolica.edu.sv/" />
<meta property="og:locale" content="es_ES" />
<meta property="og:type" content="website" />
<meta property="og:title" content="Universidad Católica de El Salvador - UNICAES" />
<meta property="og:description" content="La UNICAES es una Institución de educación superior que forma profesionales integrales, con principios cristianos y conocimientos técnicos y científicos" />
<meta property="og:url" content="http://www.catolica.edu.sv/" />
<meta property="og:site_name" content="UNICAES" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras-300x269.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cca.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/LOGO-AUPRIDES-v11-300x274.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype1.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-ODUCAL-Fondo-Transparente1-300x80.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Catholic-Higher-Education.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-HACU-144x300.gif" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_UPAEP-300x78.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/AmityInstitute.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-vector-universidad-navarra-300x152.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/neiu_wordmark_color-300x51.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg-150x150.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-150x150.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-300x61.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-300x74.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-300x130.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen-300x150.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices-1-300x248.jpg" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/ccaa-300x252.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype-300x264.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro-300x199.png" />
<meta property="og:image" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-300x300.png" />
<meta name="twitter:card" content="summary" />
<meta name="twitter:description" content="La UNICAES es una Institución de educación superior que forma profesionales integrales, con principios cristianos y conocimientos técnicos y científicos" />
<meta name="twitter:title" content="Universidad Católica de El Salvador - UNICAES" />
<meta name="twitter:image" content="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" />
<script type='application/ld+json'>{"@context":"http:\/\/schema.org","@type":"WebSite","@id":"#website","url":"http:\/\/www.catolica.edu.sv\/","name":"UNICAES","potentialAction":{"@type":"SearchAction","target":"http:\/\/www.catolica.edu.sv\/?s={search_term_string}","query-input":"required name=search_term_string"}}</script>
<script type='application/ld+json'>{"@context":"http:\/\/schema.org","@type":"Organization","url":"http:\/\/www.catolica.edu.sv\/","sameAs":["https:\/\/www.facebook.com\/UNICAES\/"],"@id":"#organization","name":"UNIVERSIDAD CATOLICA DE EL SALVADOR","logo":"http:\/\/www.catolica.edu.sv\/wp-content\/uploads\/2017\/04\/logo-UNICAES-png.png"}</script>
<!-- / Yoast SEO Premium plugin. -->

<link rel='dns-prefetch' href='//fonts.googleapis.com' />
<link rel='dns-prefetch' href='//s.w.org' />
<link rel="alternate" type="application/rss+xml" title="UNICAES &raquo; Feed" href="http://www.catolica.edu.sv/?feed=rss2" />
<link rel="alternate" type="application/rss+xml" title="UNICAES &raquo; RSS de los comentarios" href="http://www.catolica.edu.sv/?feed=comments-rss2" />
<link rel="alternate" type="text/calendar" title="UNICAES &raquo; iCal Feed" href="http://www.catolica.edu.sv?post_type=tribe_events&#038;ical=1" />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.2.1\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/www.catolica.edu.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.7.9"}};
			!function(a,b,c){function d(a){var b,c,d,e,f=String.fromCharCode;if(!k||!k.fillText)return!1;switch(k.clearRect(0,0,j.width,j.height),k.textBaseline="top",k.font="600 32px Arial",a){case"flag":return k.fillText(f(55356,56826,55356,56819),0,0),!(j.toDataURL().length<3e3)&&(k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,65039,8205,55356,57096),0,0),b=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55356,57331,55356,57096),0,0),c=j.toDataURL(),b!==c);case"emoji4":return k.fillText(f(55357,56425,55356,57341,8205,55357,56507),0,0),d=j.toDataURL(),k.clearRect(0,0,j.width,j.height),k.fillText(f(55357,56425,55356,57341,55357,56507),0,0),e=j.toDataURL(),d!==e}return!1}function e(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var f,g,h,i,j=b.createElement("canvas"),k=j.getContext&&j.getContext("2d");for(i=Array("flag","emoji4"),c.supports={everything:!0,everythingExceptFlag:!0},h=0;h<i.length;h++)c.supports[i[h]]=d(i[h]),c.supports.everything=c.supports.everything&&c.supports[i[h]],"flag"!==i[h]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[i[h]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(g=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",g,!1),a.addEventListener("load",g,!1)):(a.attachEvent("onload",g),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),f=c.source||{},f.concatemoji?e(f.concatemoji):f.wpemoji&&f.twemoji&&(e(f.twemoji),e(f.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='stylesheet' id='contact-form-7-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/contact-form-7/includes/css/styles.css?ver=4.7' type='text/css' media='all' />
<link rel='stylesheet' id='rs-plugin-settings-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/css/settings.css?ver=5.2.5' type='text/css' media='all' />
<style id='rs-plugin-settings-inline-css' type='text/css'>
#rs-demo-id {}
</style>
<link rel='stylesheet' id='tribe-events-calendar-style-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/the-events-calendar/src/resources/css/tribe-events-full.min.css?ver=4.6.10.1' type='text/css' media='all' />
<link rel='stylesheet' id='tribe-events-calendar-mobile-style-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/the-events-calendar/src/resources/css/tribe-events-full-mobile.min.css?ver=4.6.10.1' type='text/css' media='only screen and (max-width: 768px)' />
<link rel='stylesheet' id='xmenu-menu-amination-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/g5plus-framework/xmenu/assets/css/amination.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='slickr-flickr-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/styles/public.css?ver=2.5.4' type='text/css' media='all' />
<link rel='stylesheet' id='slickr-flickr-lightbox-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/styles/lightGallery.css?ver=1.0' type='text/css' media='all' />
<link rel='stylesheet' id='dashicons-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-includes/css/dashicons.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='thickbox-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-includes/js/thickbox/thickbox.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='galleria-classic-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/galleria/themes/classic/galleria.classic.css?ver=1.4.2' type='text/css' media='all' />
<link rel='stylesheet' id='js_composer_front-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/css/js_composer.min.css?ver=4.11.2.1' type='text/css' media='all' />
<link rel='stylesheet' id='font-awesome-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/font-awesome/css/font-awesome.min.css?ver=4.11.2.1' type='text/css' media='all' />
<link rel='stylesheet' id='font-awesome-animation-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/fonts-awesome/css/font-awesome-animation.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='bootstrap-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/bootstrap/css/bootstrap.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='owl-carousel-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/owl-carousel/assets/owl.carousel.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='prettyPhoto-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/prettyPhoto/css/prettyPhoto.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='peffect-scrollbar-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/perfect-scrollbar/css/perfect-scrollbar.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='slick-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/slick/css/slick.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='g5plus_framework_style-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/style.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='g5plus_framework_rtl-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/css/rtl.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='redux-google-fonts-g5plus_academia_options-css'  property='stylesheet' href='http://fonts.googleapis.com/css?family=Oswald%3A300%2C400%2C700&#038;ver=1510765625' type='text/css' media='all' />
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-includes/js/jquery/jquery.js?ver=1.12.4'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-includes/js/jquery/jquery-migrate.min.js?ver=1.4.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/js/jquery.themepunch.tools.min.js?ver=5.2.5'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/js/jquery.themepunch.revolution.min.js?ver=5.2.5'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/scripts/lightGallery.min.js?ver=1.0'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var thickboxL10n = {"next":"Siguiente >","prev":"< Anterior","image":"Imagen","of":"de","close":"Cerrar","noiframes":"Esta funci\u00f3n requiere de frames insertados. Tienes los iframes desactivados o tu navegador no los soporta.","loadingAnimation":"http:\/\/www.catolica.edu.sv\/wp-includes\/js\/thickbox\/loadingAnimation.gif"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-includes/js/thickbox/thickbox.js?ver=3.1-20121105'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/galleria/galleria-1.4.2.min.js?ver=1.4.2'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/galleria/themes/classic/galleria.classic.min.js?ver=1.4.2'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/scripts/responsiveslides.min.js?ver=1.54'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/slickr-flickr/scripts/public.js?ver=2.5.4'></script>
<link rel='https://api.w.org/' href='http://www.catolica.edu.sv/?rest_route=/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://www.catolica.edu.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://www.catolica.edu.sv/wp-includes/wlwmanifest.xml" /> 
<meta name="generator" content="WordPress 4.7.9" />
<link rel='shortlink' href='http://www.catolica.edu.sv/' />
<link rel="alternate" type="application/json+oembed" href="http://www.catolica.edu.sv/?rest_route=%2Foembed%2F1.0%2Fembed&#038;url=http%3A%2F%2Fwww.catolica.edu.sv%2F" />
<link rel="alternate" type="text/xml+oembed" href="http://www.catolica.edu.sv/?rest_route=%2Foembed%2F1.0%2Fembed&#038;url=http%3A%2F%2Fwww.catolica.edu.sv%2F&#038;format=xml" />
<meta name="tec-api-version" content="v1"><meta name="tec-api-origin" content="http://www.catolica.edu.sv"><link rel="https://theeventscalendar.com/" href="http://www.catolica.edu.sv/?rest_route=/tribe/events/v1/" /><style id="g5plus_custom_style" type="text/css"></style><style type="text/css">
                                     </style><meta name="generator" content="Powered by Visual Composer - drag and drop page builder for WordPress."/>
<!--[if lte IE 9]><link rel="stylesheet" type="text/css" href="http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/css/vc_lte_ie9.min.css" media="screen"><![endif]--><!--[if IE  8]><link rel="stylesheet" type="text/css" href="http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/css/vc-ie8.min.css" media="screen"><![endif]--><style type="text/css">.broken_link, a.broken_link {
	text-decoration: line-through;
}</style><meta name="generator" content="Powered by Slider Revolution 5.2.5 - responsive, Mobile-Friendly Slider Plugin for WordPress with comfortable drag and drop interface." />
<link rel="icon" href="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logoth-150x150.jpg" sizes="32x32" />
<link rel="icon" href="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logoth.jpg" sizes="192x192" />
<link rel="apple-touch-icon-precomposed" href="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logoth.jpg" />
<meta name="msapplication-TileImage" content="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logoth.jpg" />
<link rel="stylesheet" type="text/css" media="all" href="http://www.catolica.edu.sv/?custom-page=header-custom-css&amp;current_page_id=321"/><style type="text/css" title="dynamic-css" class="options-output">body{background-repeat:no-repeat;background-size:cover;background-attachment:fixed;background-position:center center;}.site-loading{background-color:;}body{font-family:Oswald;line-height:36px;font-weight:400;font-style:normal;font-size:15px;}h1{font-family:Oswald;line-height:42px;font-weight:700;font-style:normal;font-size:36px;}h2{font-family:Oswald;line-height:36px;font-weight:700;font-style:normal;font-size:27px;}h3{font-family:Oswald;line-height:29px;font-weight:400;font-style:normal;font-size:22px;}h4{font-family:Oswald;line-height:23px;font-weight:400;font-style:normal;font-size:17px;}h5{font-family:Oswald;line-height:17px;font-weight:400;font-style:normal;font-size:13px;}h6{font-family:Oswald;line-height:15px;font-weight:400;font-style:normal;font-size:11px;}{font-family:Oswald;}{font-family:Oswald;}{font-family:Oswald;}</style><style type="text/css" data-type="vc_shortcodes-custom-css">.vc_custom_1518622494109{margin-top: 0px !important;}</style><noscript><style type="text/css"> .wpb_animate_when_almost_visible { opacity: 1; }</style></noscript> 



<script>
!function(f,b,e,v,n,t,s)
{if(f.fbq)return;n=f.fbq=function(){n.callMethod?
n.callMethod.apply(n,arguments):n.queue.push(arguments)};
if(!f._fbq)f._fbq=n;n.push=n;n.loaded=!0;n.version='2.0';
n.queue=[];t=b.createElement(e);t.async=!0;
t.src=v;s=b.getElementsByTagName(e)[0];
s.parentNode.insertBefore(t,s)}(window,document,'script',
'https://connect.facebook.net/en_US/fbevents.js');
 fbq('init', '608600756196474'); 
fbq('track', 'PageView');
</script>
<noscript>
 <img height="1" width="1" 
src="https://www.facebook.com/tr?id=608600756196474&ev=PageView
&noscript=1"/>
</noscript>





	</head>
	<!-- Close Head -->
	<body class="home page-template-default page page-id-321 tribe-no-js tribe-bar-is-disabled page-loading footer-static boxed header-3 unknown wpb-js-composer js-comp-ver-4.11.2.1 vc_responsive" data-responsive="991" data-header="header-3">

		<div class="site-loading">
    <div class="block-center">
        <div class="block-center-inner">
            
                
                
                
                
                
                
                
                                    <div class="sk-fading-circle">
                        <div class="sk-circle1 sk-circle"></div>
                        <div class="sk-circle2 sk-circle"></div>
                        <div class="sk-circle3 sk-circle"></div>
                        <div class="sk-circle4 sk-circle"></div>
                        <div class="sk-circle5 sk-circle"></div>
                        <div class="sk-circle6 sk-circle"></div>
                        <div class="sk-circle7 sk-circle"></div>
                        <div class="sk-circle8 sk-circle"></div>
                        <div class="sk-circle9 sk-circle"></div>
                        <div class="sk-circle10 sk-circle"></div>
                        <div class="sk-circle11 sk-circle"></div>
                        <div class="sk-circle12 sk-circle"></div>
                    </div>
                
                        </div>
    </div>
</div>


		<!-- Open Wrapper -->
		<div id="wrapper">

		<header id="main-header-wrapper" class="main-header">
	
	<div class="header-nav-wrapper header-3">
	<div class="container">
		<div class="header-container clearfix">
			<div class="header-logo">
	<a href="http://www.catolica.edu.sv/" title="UNICAES - Universidad Católica de El Salvador">
		<img class="has-retina" style="height:50px" src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/fonlogo.jpg" alt="UNICAES - Universidad Católica de El Salvador" />
					<img class="retina-logo" style="height:50px" src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/fonlogo.jpg" alt="UNICAES - Universidad Católica de El Salvador"/>
			</a>
</div>
			<div class="header-nav-right">
									<div id="primary-menu" class="menu-wrapper">
						<ul id="main-menu" class="main-menu sub-menu-light x-nav-menu x-nav-menu_main-menu x-animate-sign-flip"><li id="menu-item-879" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-home current-menu-item page_item page-item-321 current_page_item x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Inicio</span></a></li><li id="menu-item-3079" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3063" class="x-menu-a-text"><span class="x-menu-text">Nosotros</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-882" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=390" class="x-menu-a-text"><span class="x-menu-text">Identidad Institucional</span></a></li><li id="menu-item-940" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=938" class="x-menu-a-text"><span class="x-menu-text">Reseña Histórica</span></a></li><li id="menu-item-881" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=395" class="x-menu-a-text"><span class="x-menu-text">Autoridades Universitarias</span></a></li></ul></li><li id="menu-item-2623" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://www.registroacademico.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Admisión</span></a></li><li id="menu-item-1061" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1057" class="x-menu-a-text"><span class="x-menu-text">Oferta Académica</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1010" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=669" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ingeniería y Arquitectura</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-8418" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=8367" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Desarrollo de Software</span></a></li><li id="menu-item-1164" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1159" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Telecomunicaciones y Redes</span></a></li><li id="menu-item-1169" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1144" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Civil</span></a></li><li id="menu-item-1167" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1153" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Industrial</span></a></li><li id="menu-item-1166" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1155" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Sistemas Informáticos</span></a></li><li id="menu-item-1165" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1157" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Agronómica</span></a></li><li id="menu-item-1163" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1161" class="x-menu-a-text"><span class="x-menu-text">Arquitectura</span></a></li></ul></li><li id="menu-item-1004" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=674" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias Empresariales</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1194" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1170" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas</span></a></li><li id="menu-item-3006" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2273" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas (Semipresencial)</span></a></li><li id="menu-item-1193" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1173" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Sistemas Informáticos Administrativos</span></a></li><li id="menu-item-1192" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1176" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Contaduría Pública</span></a></li><li id="menu-item-1191" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1179" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Mercadeo y Negocios Internacionales</span></a></li><li id="menu-item-1190" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1182" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Gestión y Desarrollo Turístico</span></a></li></ul></li><li id="menu-item-1009" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=676" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias y Humanidades</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1096" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1067" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Diseño Gráfico Publicitario</span></a></li><li id="menu-item-1097" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1065" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias Jurídicas</span></a></li><li id="menu-item-1095" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1069" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Periodismo y Comunicación Audiovisual</span></a></li><li id="menu-item-1094" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1071" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias Religiosas</span></a></li><li id="menu-item-1092" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1075" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Idioma Inglés</span></a></li><li id="menu-item-1090" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1079" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés</span></a></li><li id="menu-item-1093" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1073" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica</span></a></li><li id="menu-item-3018" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3011" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés (Semipresencial)</span></a></li><li id="menu-item-3024" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3021" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica (Semipresencial)</span></a></li><li id="menu-item-1091" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1077" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Matemática (Semipresencial)</span></a></li><li id="menu-item-1089" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1081" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Dirección y Administración Escolar (Semipresencial)</span></a></li></ul></li><li id="menu-item-1008" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=667" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias de la Salud</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1143" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1132" class="x-menu-a-text"><span class="x-menu-text">Doctorado en Medicina</span></a></li><li id="menu-item-1142" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1137" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Enfermería</span></a></li><li id="menu-item-1141" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1139" class="x-menu-a-text"><span class="x-menu-text">Técnico en Enfermería</span></a></li></ul></li><li id="menu-item-3042" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3028" class="x-menu-a-text"><span class="x-menu-text">Carreras semipresenciales</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-3056" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3054" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés (semipresencial)</span></a></li><li id="menu-item-3046" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3043" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas (semipresencial)</span></a></li><li id="menu-item-3051" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3047" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica (semipresencial)</span></a></li><li id="menu-item-3053" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3050" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Dirección y Administración Escolar (semipresencial)</span></a></li><li id="menu-item-3060" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3057" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Matemática (semipresencial)</span></a></li></ul></li></ul></li><li id="menu-item-999" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=671" class="x-menu-a-text"><span class="x-menu-text">Maestrías</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1480" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1446" class="x-menu-a-text"><span class="x-menu-text">Maestría en Asesoría Educativa</span></a></li><li id="menu-item-1479" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1449" class="x-menu-a-text"><span class="x-menu-text">Maestría en Dirección Estratégica de Empresas</span></a></li><li id="menu-item-1482" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1432" class="x-menu-a-text"><span class="x-menu-text">Maestría en Gestión y Desarrollo Turístico</span></a></li><li id="menu-item-1481" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1438" class="x-menu-a-text"><span class="x-menu-text">Maestría en Gerencia y Gestión Ambiental</span></a></li><li id="menu-item-9170" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=9092" class="x-menu-a-text"><span class="x-menu-text">Becas Maestrías</span></a></li><li id="menu-item-1771" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1737" class="x-menu-a-text"><span class="x-menu-text">Diplomados y Cursos</span></a></li></ul></li><li id="menu-item-1023" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1017" class="x-menu-a-text"><span class="x-menu-text">Unidades</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-2622" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://www.bibliotecaunicaes.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Biblioteca Miguel de Cervantes</span></a></li><li id="menu-item-1026" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1024" class="x-menu-a-text"><span class="x-menu-text">Departamento de Idiomas</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-1040" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1038" class="x-menu-a-text"><span class="x-menu-text">Inglés</span></a></li><li id="menu-item-2617" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2612" class="x-menu-a-text"><span class="x-menu-text">Francés</span></a></li><li id="menu-item-2616" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2614" class="x-menu-a-text"><span class="x-menu-text">Mandarín</span></a></li></ul></li><li id="menu-item-981" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a target="_blank" href="http://www.diyps.catolica.edu.sv" class="x-menu-a-text"><span class="x-menu-text">Dirección de Investigación y Proyección Social</span></a></li><li id="menu-item-2644" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2639" class="x-menu-a-text"><span class="x-menu-text">Evaluación y Currículo</span></a></li><li id="menu-item-3210" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3201" class="x-menu-a-text"><span class="x-menu-text">American Space</span></a></li><li id="menu-item-6346" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://registroacademico.catolica.edu.sv" class="x-menu-a-text"><span class="x-menu-text">Registro Académico</span></a></li><li id="menu-item-2762" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1368" class="x-menu-a-text"><span class="x-menu-text">Bienestar Universitario</span></a></li><li id="menu-item-2233" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2231" class="x-menu-a-text"><span class="x-menu-text">Centro de Orientación de Carreras</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-6023" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=5994" class="x-menu-a-text"><span class="x-menu-text">Oportunidades de Empleo y Pasantías</span></a></li></ul></li><li id="menu-item-2235" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2227" class="x-menu-a-text"><span class="x-menu-text">Clínica Universitaria</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-9344" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=9312" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Bioquímica</span></a></li></ul></li><li id="menu-item-2643" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2641" class="x-menu-a-text"><span class="x-menu-text">Colegio Madre de la Iglesia</span></a></li><li id="menu-item-4483" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=4478" class="x-menu-a-text"><span class="x-menu-text">Colecturía</span></a></li><li id="menu-item-1472" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1407" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Tecnología Informática</span></a></li><li id="menu-item-1473" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1405" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Tejidos y Cultivos</span></a></li><li id="menu-item-1466" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1411" class="x-menu-a-text"><span class="x-menu-text">Oficina de Asesoría Legal Católica (OFALCA)</span></a></li><li id="menu-item-1468" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1419" class="x-menu-a-text"><span class="x-menu-text">Parroquia Universitaria</span></a></li><li id="menu-item-1469" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1409" class="x-menu-a-text"><span class="x-menu-text">Unidad de Comunicaciones y Mercadeo</span></a></li><li id="menu-item-1474" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1415" class="x-menu-a-text"><span class="x-menu-text">Librería UNICAES</span></a></li><li id="menu-item-2234" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2229" class="x-menu-a-text"><span class="x-menu-text">Unidad de Servicios Generales</span></a></li><li id="menu-item-1467" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1413" class="x-menu-a-text"><span class="x-menu-text">Oficina de Asesoría Psicológica y Educativa</span></a></li></ul></li><li id="menu-item-2169" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=861" class="x-menu-a-text"><span class="x-menu-text">Noticias</span></a></li><li id="menu-item-892" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=738" class="x-menu-a-text"><span class="x-menu-text">Contáctanos</span></a></li></ul>					</div>
									<div class="header-customize header-customize-nav">
		<div class="search-button-wrapper header-customize-item style-">
	<a class="icon-search-menu" href="#" data-search-type="standard"><i class="fa fa-search"></i></a>
</div><div class="header-customize-item header-social-profile-wrapper">
	<ul>
		<li><a href="https://twitter.com/unicaes_sv/" target="_blank"><i class="fa fa-twitter"></i></a></li>
<li><a href="https://www.facebook.com/UNICAES/" target="_blank"><i class="fa fa-facebook"></i></a></li>
<li><a href="https://www.youtube.com/channel/UCXDsbngj7qUa2wVlm9ogPvw" target="_blank"><i class="fa fa-youtube"></i></a></li>
<li><a href="https://www.instagram.com/UNICAES_SV/" target="_blank"><i class="fa fa-instagram"></i></a></li>
	</ul>
</div>
	</div>
			</div>
		</div>
	</div>
</div>			<div class="top-bar">
	<div class="container">
		<div class="row">
										<div class="sidebar top-bar-right col-md-12">
					<aside id="text-8" class="widget widget_text">			<div class="textwidget"><div style="color: #FFF; margin-left: -480px; position:absolute">
<h2>Universidad Católica de El Salvador</h2>

</div>
<ul class="top-bar-info">
	<li><a href="mailto:catolica@catolica.edu.sv"><i class="fa fa-paper-plane"></i> catolica@catolica.edu.sv</a></li>
	<li><i class="fa fa-clock-o"></i> Lunes - Viernes: 8:00 a.m. - 6:00 p.m. Sábado: 8:00 a.m. - 12:00 p.m.</li>
</ul></div>
		</aside>				</div>
					</div>
	</div>
</div>	</header><header id="mobile-header-wrapper" class="mobile-header header-mobile-1">
		<div class="header-container-wrapper header-mobile-sticky">
	<div class="container header-mobile-container">
		<div class="header-mobile-inner">
			<div class="toggle-icon-wrapper toggle-mobile-menu" data-ref="nav-menu-mobile" data-drop-type="fly">
				<div class="toggle-icon"> <span></span></div>
			</div>
			<div class="header-customize">
									<div class="search-button-wrapper header-customize-item">
	<a class="icon-search-menu" href="#" data-search-type="standard"><i class="fa fa-search"></i></a>
</div>											</div>
			<div class="header-logo-mobile">
	<a href="http://www.catolica.edu.sv/" title="UNICAES - Universidad Católica de El Salvador">
		<img class="has-retina" style="height:70px" src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/UNICAES_New_Logo_08.jpg" alt="UNICAES - Universidad Católica de El Salvador" />
					<img class="retina-logo" style="height:70px" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logoth.jpg" alt="UNICAES - Universidad Católica de El Salvador" />
			</a>
</div>		</div>
		<div id="nav-menu-mobile" class="header-mobile-nav menu-drop-fly">
			<form class="search-form-menu-mobile"  method="get" action="http://www.catolica.edu.sv/">
			<input type="text" name="s" placeholder="Search...">
			<button type="submit"><i class="fa fa-search"></i></button>
		</form>
					<ul id="menu-main-menu" class="nav-menu-mobile x-nav-menu x-nav-menu_main-menu x-animate-sign-flip"><li id="menu-item-mobile-879" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-home current-menu-item page_item page-item-321 current_page_item x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Inicio</span></a></li><li id="menu-item-mobile-3079" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3063" class="x-menu-a-text"><span class="x-menu-text">Nosotros</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-882" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=390" class="x-menu-a-text"><span class="x-menu-text">Identidad Institucional</span></a></li><li id="menu-item-mobile-940" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=938" class="x-menu-a-text"><span class="x-menu-text">Reseña Histórica</span></a></li><li id="menu-item-mobile-881" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=395" class="x-menu-a-text"><span class="x-menu-text">Autoridades Universitarias</span></a></li></ul></li><li id="menu-item-mobile-2623" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://www.registroacademico.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Admisión</span></a></li><li id="menu-item-mobile-1061" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1057" class="x-menu-a-text"><span class="x-menu-text">Oferta Académica</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1010" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=669" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ingeniería y Arquitectura</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-8418" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=8367" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Desarrollo de Software</span></a></li><li id="menu-item-mobile-1164" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1159" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Telecomunicaciones y Redes</span></a></li><li id="menu-item-mobile-1169" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1144" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Civil</span></a></li><li id="menu-item-mobile-1167" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1153" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Industrial</span></a></li><li id="menu-item-mobile-1166" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1155" class="x-menu-a-text"><span class="x-menu-text">Ingeniería en Sistemas Informáticos</span></a></li><li id="menu-item-mobile-1165" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1157" class="x-menu-a-text"><span class="x-menu-text">Ingeniería Agronómica</span></a></li><li id="menu-item-mobile-1163" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1161" class="x-menu-a-text"><span class="x-menu-text">Arquitectura</span></a></li></ul></li><li id="menu-item-mobile-1004" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=674" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias Empresariales</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1194" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1170" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas</span></a></li><li id="menu-item-mobile-3006" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2273" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas (Semipresencial)</span></a></li><li id="menu-item-mobile-1193" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1173" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Sistemas Informáticos Administrativos</span></a></li><li id="menu-item-mobile-1192" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1176" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Contaduría Pública</span></a></li><li id="menu-item-mobile-1191" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1179" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Mercadeo y Negocios Internacionales</span></a></li><li id="menu-item-mobile-1190" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1182" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Gestión y Desarrollo Turístico</span></a></li></ul></li><li id="menu-item-mobile-1009" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=676" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias y Humanidades</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1096" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1067" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Diseño Gráfico Publicitario</span></a></li><li id="menu-item-mobile-1097" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1065" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias Jurídicas</span></a></li><li id="menu-item-mobile-1095" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1069" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Periodismo y Comunicación Audiovisual</span></a></li><li id="menu-item-mobile-1094" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1071" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias Religiosas</span></a></li><li id="menu-item-mobile-1092" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1075" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Idioma Inglés</span></a></li><li id="menu-item-mobile-1090" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1079" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés</span></a></li><li id="menu-item-mobile-1093" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1073" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica</span></a></li><li id="menu-item-mobile-3018" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3011" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés (Semipresencial)</span></a></li><li id="menu-item-mobile-3024" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3021" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica (Semipresencial)</span></a></li><li id="menu-item-mobile-1091" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1077" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Matemática (Semipresencial)</span></a></li><li id="menu-item-mobile-1089" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1081" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Dirección y Administración Escolar (Semipresencial)</span></a></li></ul></li><li id="menu-item-mobile-1008" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=667" class="x-menu-a-text"><span class="x-menu-text">Facultad de Ciencias de la Salud</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1143" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1132" class="x-menu-a-text"><span class="x-menu-text">Doctorado en Medicina</span></a></li><li id="menu-item-mobile-1142" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1137" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Enfermería</span></a></li><li id="menu-item-mobile-1141" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1139" class="x-menu-a-text"><span class="x-menu-text">Técnico en Enfermería</span></a></li></ul></li><li id="menu-item-mobile-3042" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3028" class="x-menu-a-text"><span class="x-menu-text">Carreras semipresenciales</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-3056" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3054" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Idioma Inglés (semipresencial)</span></a></li><li id="menu-item-mobile-3046" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3043" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Administración de Empresas (semipresencial)</span></a></li><li id="menu-item-mobile-3051" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3047" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Educación Básica (semipresencial)</span></a></li><li id="menu-item-mobile-3053" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3050" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Dirección y Administración Escolar (semipresencial)</span></a></li><li id="menu-item-mobile-3060" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3057" class="x-menu-a-text"><span class="x-menu-text">Licenciatura en Ciencias de la Educación con Especialidad en Matemática (semipresencial)</span></a></li></ul></li></ul></li><li id="menu-item-mobile-999" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=671" class="x-menu-a-text"><span class="x-menu-text">Maestrías</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1480" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1446" class="x-menu-a-text"><span class="x-menu-text">Maestría en Asesoría Educativa</span></a></li><li id="menu-item-mobile-1479" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1449" class="x-menu-a-text"><span class="x-menu-text">Maestría en Dirección Estratégica de Empresas</span></a></li><li id="menu-item-mobile-1482" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1432" class="x-menu-a-text"><span class="x-menu-text">Maestría en Gestión y Desarrollo Turístico</span></a></li><li id="menu-item-mobile-1481" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1438" class="x-menu-a-text"><span class="x-menu-text">Maestría en Gerencia y Gestión Ambiental</span></a></li><li id="menu-item-mobile-9170" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=9092" class="x-menu-a-text"><span class="x-menu-text">Becas Maestrías</span></a></li><li id="menu-item-mobile-1771" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1737" class="x-menu-a-text"><span class="x-menu-text">Diplomados y Cursos</span></a></li></ul></li><li id="menu-item-mobile-1023" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1017" class="x-menu-a-text"><span class="x-menu-text">Unidades</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-2622" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://www.bibliotecaunicaes.catolica.edu.sv/" class="x-menu-a-text"><span class="x-menu-text">Biblioteca Miguel de Cervantes</span></a></li><li id="menu-item-mobile-1026" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1024" class="x-menu-a-text"><span class="x-menu-text">Departamento de Idiomas</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-1040" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1038" class="x-menu-a-text"><span class="x-menu-text">Inglés</span></a></li><li id="menu-item-mobile-2617" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2612" class="x-menu-a-text"><span class="x-menu-text">Francés</span></a></li><li id="menu-item-mobile-2616" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2614" class="x-menu-a-text"><span class="x-menu-text">Mandarín</span></a></li></ul></li><li id="menu-item-mobile-981" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a target="_blank" href="http://www.diyps.catolica.edu.sv" class="x-menu-a-text"><span class="x-menu-text">Dirección de Investigación y Proyección Social</span></a></li><li id="menu-item-mobile-2644" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2639" class="x-menu-a-text"><span class="x-menu-text">Evaluación y Currículo</span></a></li><li id="menu-item-mobile-3210" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=3201" class="x-menu-a-text"><span class="x-menu-text">American Space</span></a></li><li id="menu-item-mobile-6346" class="menu-item menu-item-type-custom menu-item-object-custom x-menu-item x-item-menu-standard"><a href="http://registroacademico.catolica.edu.sv" class="x-menu-a-text"><span class="x-menu-text">Registro Académico</span></a></li><li id="menu-item-mobile-2762" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1368" class="x-menu-a-text"><span class="x-menu-text">Bienestar Universitario</span></a></li><li id="menu-item-mobile-2233" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2231" class="x-menu-a-text"><span class="x-menu-text">Centro de Orientación de Carreras</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-6023" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=5994" class="x-menu-a-text"><span class="x-menu-text">Oportunidades de Empleo y Pasantías</span></a></li></ul></li><li id="menu-item-mobile-2235" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-has-children x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2227" class="x-menu-a-text"><span class="x-menu-text">Clínica Universitaria</span><b class="x-caret"></b></a>			<ul class="x-sub-menu x-sub-menu-standard x-list-style-none">
		<li id="menu-item-mobile-9344" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=9312" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Bioquímica</span></a></li></ul></li><li id="menu-item-mobile-2643" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2641" class="x-menu-a-text"><span class="x-menu-text">Colegio Madre de la Iglesia</span></a></li><li id="menu-item-mobile-4483" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=4478" class="x-menu-a-text"><span class="x-menu-text">Colecturía</span></a></li><li id="menu-item-mobile-1472" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1407" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Tecnología Informática</span></a></li><li id="menu-item-mobile-1473" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1405" class="x-menu-a-text"><span class="x-menu-text">Laboratorio de Tejidos y Cultivos</span></a></li><li id="menu-item-mobile-1466" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1411" class="x-menu-a-text"><span class="x-menu-text">Oficina de Asesoría Legal Católica (OFALCA)</span></a></li><li id="menu-item-mobile-1468" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1419" class="x-menu-a-text"><span class="x-menu-text">Parroquia Universitaria</span></a></li><li id="menu-item-mobile-1469" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1409" class="x-menu-a-text"><span class="x-menu-text">Unidad de Comunicaciones y Mercadeo</span></a></li><li id="menu-item-mobile-1474" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1415" class="x-menu-a-text"><span class="x-menu-text">Librería UNICAES</span></a></li><li id="menu-item-mobile-2234" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=2229" class="x-menu-a-text"><span class="x-menu-text">Unidad de Servicios Generales</span></a></li><li id="menu-item-mobile-1467" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=1413" class="x-menu-a-text"><span class="x-menu-text">Oficina de Asesoría Psicológica y Educativa</span></a></li></ul></li><li id="menu-item-mobile-2169" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=861" class="x-menu-a-text"><span class="x-menu-text">Noticias</span></a></li><li id="menu-item-mobile-892" class="menu-item menu-item-type-post_type menu-item-object-page x-menu-item x-item-menu-standard"><a href="http://www.catolica.edu.sv/?page_id=738" class="x-menu-a-text"><span class="x-menu-text">Contáctanos</span></a></li></ul>	
	</div>
	<div class="main-menu-overlay"></div>
	</div>
</div></header>	<div id="search_popup_wrapper" class="dialog">
		<div class="dialog__overlay"></div>
		<div class="dialog__content">
			<div class="morph-shape">
				<svg xmlns="http://www.w3.org/2000/svg" width="100%" height="100%" viewBox="0 0 520 280"
				     preserveAspectRatio="none">
					<rect x="3" y="3" fill="none" width="516" height="276"/>
				</svg>
			</div>
			<div class="dialog-inner">
				<h2>Enter your keyword</h2>
				<form  method="get" action="http://www.catolica.edu.sv/" class="search-popup-inner">
					<input type="text" name="s" placeholder="Search...">
					<button type="submit">Search</button>
				</form>
				<div><button class="action" data-dialog-close="close" type="button"><i class="fa fa-close"></i></button></div>
			</div>
		</div>
	</div>

			<!-- Open Wrapper Content -->
			<div id="wrapper-content" class="clearfix">

			<main  class="site-content-page">
									<div class="site-content-page-inner ">
				<div class="page-content">
                    <div id="post-321" class="post-321 page type-page status-publish hentry">
	<div class="entry-content clearfix">
		<div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12 vc_hidden-sm vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="wpb_revslider_element wpb_content_element"><link href="http://fonts.googleapis.com/css?family=Roboto%3A500" rel="stylesheet" property="stylesheet" type="text/css" media="all" /><link href="http://fonts.googleapis.com/css?family=Oswald%3A400%2C500%2C300%2C900" rel="stylesheet" property="stylesheet" type="text/css" media="all" />
<div id="rev_slider_3_1_wrapper" class="rev_slider_wrapper fullwidthbanner-container" style="margin:0px auto;background-color:transparent;padding:0px;margin-top:0px;margin-bottom:0px;">
<!-- START REVOLUTION SLIDER 5.2.5 auto mode -->
	<div id="rev_slider_3_1" class="rev_slider fullwidthabanner" style="display:none;" data-version="5.2.5">
<ul>	<!-- SLIDE  -->
	<li data-index="rs-68" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2018/02/Slide-Web1-100x50.png"  data-delay="8000"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/Slide-Web1.png"  alt="" title="Slide Web(1)"  width="1200" height="700" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption aca rev-btn " 
			 id="slide-68-layer-1" 
			 data-x="['left','left','left','left']" data-hoffset="['443','443','443','443']" 
			 data-y="['top','top','top','top']" data-voffset="['288','288','288','288']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(255, 255, 255, 10.00);bg:rgba(136, 12, 10, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_blank","url":"https:\/\/www.moralurbanidadycivica.com\/"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			
			style="z-index: 5; white-space: nowrap; font-size: 25px; line-height: 20px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:Roboto;background-color:rgba(0, 0, 0, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);border-radius:3px 3px 3px 3px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">AQUÍ </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-53" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2018/01/slider-web-100x50.jpg"  data-delay="8410.000610351562"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2018/01/slider-web.jpg"  alt="" title="slider-web"  width="1200" height="700" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-53-layer-1" 
			 data-x="['left','left','left','left']" data-hoffset="['478','478','478','478']" 
			 data-y="['top','top','top','top']" data-voffset="['335','335','335','335']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			
			style="z-index: 5; white-space: nowrap; font-size: 50px;">Información de Graduación LX </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption rev-btn rev-withicon " 
			 id="slide-53-layer-2" 
			 data-x="['left','left','left','left']" data-hoffset="['698','698','698','698']" 
			 data-y="['top','top','top','top']" data-voffset="['417','417','417','417']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":" http:\/\/www.catolica.edu.sv\/?tribe_events=informacion-graduacion-lx"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			
			style="z-index: 6; white-space: nowrap; font-size: 45px; line-height: 17px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:oswald;background-color:rgba(136, 12, 10, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);border-radius:30px 30px 30px 30px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">Aquí<i class="fa-icon-chevron-right"></i> </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-8" data-transition="curtain-2,boxslide,slidedown" data-slotamount="default,default,default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default,default,default" data-easeout="default,default,default" data-masterspeed="default,default,default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/07/web1-100x50.png"  data-delay="8130"  data-rotate="0,0,0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/07/web1.png"  alt="" title="web1"  width="1200" height="700" data-bgposition="center bottom" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-sub-heading-top   tp-resizeme" 
			 id="slide-8-layer-2" 
			 data-x="['left','center','center','center']" data-hoffset="['652','84','-30','-117']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-252','-264','-265','-273']" 
						data-fontsize="['30','28','28','28']"
			data-width="['262','none','none','none']"
			data-height="['65','none','none','none']"
			data-whitespace="['normal','nowrap','nowrap','nowrap']"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="649.6875" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.6875" 

			style="z-index: 5; min-width: 262px; max-width: 262px; max-width: 65px; max-width: 65px; white-space: normal; font-size: 30px; color: rgba(49, 52, 73, 1.00);">CONOCE NUESTRO </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-8-layer-1" 
			 data-x="['left','center','center','center']" data-hoffset="['651','232','81','24']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-229','-222','-228','-238']" 
						data-fontsize="['50','60','50','45']"
			data-lineheight="['72','72','72','54']"
			data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="899.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 6; white-space: nowrap; font-size: 50px; color: rgba(49, 52, 73, 1.00);">CAMPUS UNICAES </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption academia-sub-heading-bottom   tp-resizeme" 
			 id="slide-8-layer-3" 
			 data-x="['left','center','center','center']" data-hoffset="['714','281','46','76']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-191','-183','-182','-206']" 
						data-color="['rgba(6, 2, 10, 1.00)','rgba(13, 0, 33, 1.00)','rgba(13, 0, 33, 1.00)','rgba(13, 0, 33, 1.00)']"
			data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="x:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;s:1500;e:Power3.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:0px;s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="1149.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 7; white-space: nowrap; color: rgba(6, 2, 10, 1.00);font-family:Oswald;">Y NUESTRAS CARRERAS UNIVERSITARIAS </div>

		<!-- LAYER NR. 4 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-8-layer-6" 
			 data-x="['left','center','center','center']" data-hoffset="['676','176','-3','-53']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-137','-132','-128','-157']" 
						data-fontsize="['16','16','16','12']"
			data-lineheight="['30','22','22','22']"
			data-fontweight="['300','400','400','400']"
			data-color="['rgba(2, 2, 2, 1.00)','rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)']"
			data-width="['141','none','none','none']"
			data-height="none"
			data-whitespace="['normal','nowrap','nowrap','nowrap']"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(255, 255, 255, 1.00);bg:rgba(136, 12, 10, 1.00);"
 
			 data-transform_in="opacity:0;s:1500;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1010;e:Power2.easeInOut;" 
			data-start="1149.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=1057"}]'
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 8; min-width: 141px; max-width: 141px; white-space: normal; font-size: 16px; line-height: 30px; font-weight: 300; color: rgba(2, 2, 2, 1.00);font-family:Oswald;text-align:center;background-color:rgba(237, 189, 63, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">PREGRADOS </div>

		<!-- LAYER NR. 5 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-8-layer-8" 
			 data-x="['left','center','center','center']" data-hoffset="['843','351','173','111']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-137','-138','-127','-159']" 
						data-fontsize="['16','16','16','12']"
			data-lineheight="['30','22','22','22']"
			data-fontweight="['300','400','400','500']"
			data-width="['141','none','none','none']"
			data-height="none"
			data-whitespace="['normal','nowrap','nowrap','nowrap']"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(10, 0, 2, 1.00);bg:rgba(237, 189, 63, 1.00);"
 
			 data-transform_in="opacity:0;s:1500;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1010;e:Power2.easeInOut;" 
			data-start="1399.6875" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=671"}]'
			data-responsive_offset="on" 

			 data-end="6989.6875" 

			style="z-index: 9; min-width: 141px; max-width: 141px; white-space: normal; font-size: 16px; line-height: 30px; font-weight: 300;font-family:Oswald;text-align:center;background-color:rgba(136, 12, 10, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">POSTGRADOS </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-21" data-transition="slidedown" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/07/web2-100x50.png"  data-delay="8220"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/07/web2.png"  alt="" title="web2"  width="1200" height="700" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption rev-btn " 
			 id="slide-21-layer-4" 
			 data-x="['left','left','left','left']" data-hoffset="['318','318','318','318']" 
			 data-y="['top','top','top','top']" data-voffset="['193','193','193','193']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?post_type=tribe_events"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			 data-end="7860" 

			style="z-index: 5; white-space: nowrap; font-size: 35px; line-height: 25px; font-weight: 500; color: rgba(12, 12, 12, 1.00);font-family:oswald;background-color:rgba(237, 189, 63, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">EVENTOS </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption rev-btn " 
			 id="slide-21-layer-5" 
			 data-x="['left','left','left','left']" data-hoffset="['572','572','572','572']" 
			 data-y="['top','top','top','top']" data-voffset="['193','193','193','193']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=861"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			 data-end="7900" 

			style="z-index: 6; white-space: nowrap; font-size: 35px; line-height: 25px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:oswald;background-color:rgba(136, 12, 10, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">NOTICIAS </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-21-layer-6" 
			 data-x="['left','left','left','left']" data-hoffset="['404','404','404','404']" 
			 data-y="['top','top','top','top']" data-voffset="['110','110','110','110']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="7870" 

			style="z-index: 7; white-space: nowrap; color: rgba(12, 12, 12, 1.00);">ENTÉRATE DE: </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-7" data-transition="curtain-1,boxfade,slidedown" data-slotamount="default,default,default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default,default,default" data-easeout="default,default,default" data-masterspeed="default,default,default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2016/07/unnamed-100x50.jpg"  data-delay="9000"  data-rotate="0,0,0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2016/07/unnamed.jpg"  alt="" title="unnamed"  width="1173" height="782" data-bgposition="right center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-7-layer-1" 
			 data-x="['left','left','left','left']" data-hoffset="['71','64','47','32']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-171','-186','-186','-235']" 
						data-fontsize="['60','60','50','30']"
			data-lineheight="['72','72','72','60']"
			data-width="['843','844','844','399']"
			data-height="['145','none','none','none']"
			data-whitespace="normal"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1000;e:Power2.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="650" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="8360" 

			style="z-index: 5; min-width: 843px; max-width: 843px; max-width: 145px; max-width: 145px; white-space: normal; color: rgba(10, 10, 10, 1.00);">CENTRO REGIONAL DE ILOBASCO </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption academia-sub-heading   tp-resizeme" 
			 id="slide-7-layer-2" 
			 data-x="['left','left','left','left']" data-hoffset="['72','63','46','31']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-260','-236','-229','-268']" 
						data-fontsize="['65','75','75','35']"
			data-width="['345','339','339','240']"
			data-height="['58','83','83','54']"
			data-whitespace="normal"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1000;e:Power2.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="900" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="8009.8965454102" 

			style="z-index: 6; min-width: 345px; max-width: 345px; max-width: 58px; max-width: 58px; white-space: normal; font-size: 65px; line-height: 50px; color: rgba(10, 10, 10, 1.00);">UNICAES </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-7-layer-4" 
			 data-x="['left','left','left','left']" data-hoffset="['398','335','286','218']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-140','-125','-129','-187']" 
						data-fontsize="['20','20','20','12']"
			data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(10, 2, 4, 1.00);bg:rgba(237, 189, 63, 1.00);"
 
			 data-transform_in="opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1000;e:Power2.easeIn;" 
			data-start="1400" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.cri.catolica.edu.sv\/"}]'
			data-responsive_offset="on" 

			 data-end="7000" 

			style="z-index: 7; white-space: nowrap; font-size: 20px;font-family:Oswald;background-color:rgba(136, 12, 10, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">Ir al sitio web </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-47" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/05/prueba2-100x50.jpg"  data-delay="10000"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/05/prueba2.jpg"  alt="" title="prueba2"  width="1200" height="700" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption rev-btn rev-hiddenicon  tp-resizeme" 
			 id="slide-47-layer-2" 
			 data-x="['center','center','center','center']" data-hoffset="['11','11','11','11']" 
			 data-y="['top','top','top','top']" data-voffset="['99','99','99','99']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);td:overline;bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=7577"}]'
			data-responsive_offset="on" 

			
			style="z-index: 5; white-space: nowrap; font-size: 55px; line-height: 20px; font-weight: 900; color: rgba(214, 240, 47, 1.00);font-family:oswald;text-align:center;text-transform:uppercase;background-color:rgba(1, 15, 90, 1.00);padding:25px 55px 25px 55px;border-color:rgba(0, 0, 0, 1.00);border-radius:30px 30px 30px 30px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;letter-spacing:1px;cursor:pointer;">Haz clic <i class="fa-icon-mouse-pointer"></i> </div>
	</li>
</ul>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss="";
						if(htmlDiv) {
							htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
						}else{
							var htmlDiv = document.createElement("div");
							htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
							document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
						}
					</script>
<div class="tp-bannertimer tp-bottom" style="visibility: hidden !important;"></div>	</div>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss=".tp-caption.academia-sub-heading-top,.academia-sub-heading-top{color:rgba(255,255,255,1.00);font-size:28px;line-height:33.6px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left}.tp-caption.academia-heading,.academia-heading{color:rgba(255,255,255,1.00);font-size:60px;line-height:72px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left;letter-spacing:0.02em}.tp-caption.academia-sub-heading-bottom,.academia-sub-heading-bottom{color:rgba(255,255,255,1.00);font-size:16px;line-height:19.2px;font-weight:400;font-style:normal;font-family:Roboto;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left}.tp-caption.academia-button-bg,.academia-button-bg{color:rgba(255,255,255,1.00);font-size:12px;line-height:22px;font-weight:400;font-style:normal;font-family:Roboto;padding:11px 30px 11px 30px;text-decoration:none;background-color:rgba(47,167,203,1.00);border-color:transparent;border-style:solid;border-width:0px;border-radius:0px 0px 0px 0px;text-align:left;letter-spacing:0.05em !important;-webkit-transition:all .3s !important;-moz-transition:all .3s !important;-o-transition:all .3s !important;transition:all .3s !important}.tp-caption.academia-button-bg:hover,.academia-button-bg:hover{color:rgba(255,255,255,1.00);text-decoration:none;background-color:rgba(145,95,169,1.00);border-color:transparent;border-style:none;border-width:0px;border-radius:0px 0px 0px 0px}.tp-caption.academia-sub-heading,.academia-sub-heading{color:rgba(255,255,255,1.00);font-size:24px;line-height:28.8px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left;letter-spacing:0.1em}";
				if(htmlDiv) {
					htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
				}else{
					var htmlDiv = document.createElement("div");
					htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
					document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
				}
			</script>
		<script type="text/javascript">
						/******************************************
				-	PREPARE PLACEHOLDER FOR SLIDER	-
			******************************************/

			var setREVStartSize=function(){
				try{var e=new Object,i=jQuery(window).width(),t=9999,r=0,n=0,l=0,f=0,s=0,h=0;
					e.c = jQuery('#rev_slider_3_1');
					e.responsiveLevels = [1240,1024,778,480];
					e.gridwidth = [1200,1024,778,480];
					e.gridheight = [700,650,600,600];
							
					e.sliderLayout = "auto";
					if(e.responsiveLevels&&(jQuery.each(e.responsiveLevels,function(e,f){f>i&&(t=r=f,l=e),i>f&&f>r&&(r=f,n=e)}),t>r&&(l=n)),f=e.gridheight[l]||e.gridheight[0]||e.gridheight,s=e.gridwidth[l]||e.gridwidth[0]||e.gridwidth,h=i/s,h=h>1?1:h,f=Math.round(h*f),"fullscreen"==e.sliderLayout){var u=(e.c.width(),jQuery(window).height());if(void 0!=e.fullScreenOffsetContainer){var c=e.fullScreenOffsetContainer.split(",");if (c) jQuery.each(c,function(e,i){u=jQuery(i).length>0?u-jQuery(i).outerHeight(!0):u}),e.fullScreenOffset.split("%").length>1&&void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0?u-=jQuery(window).height()*parseInt(e.fullScreenOffset,0)/100:void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0&&(u-=parseInt(e.fullScreenOffset,0))}f=u}else void 0!=e.minHeight&&f<e.minHeight&&(f=e.minHeight);e.c.closest(".rev_slider_wrapper").css({height:f})
					
				}catch(d){console.log("Failure at Presize of Slider:"+d)}
			};
			
			setREVStartSize();
			
						var tpj=jQuery;
			
			var revapi3;
			tpj(document).ready(function() {
				if(tpj("#rev_slider_3_1").revolution == undefined){
					revslider_showDoubleJqueryError("#rev_slider_3_1");
				}else{
					revapi3 = tpj("#rev_slider_3_1").show().revolution({
						sliderType:"standard",
jsFileLocation:"//www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/js/",
						sliderLayout:"auto",
						dottedOverlay:"none",
						delay:4000,
						navigation: {
							keyboardNavigation:"off",
							keyboard_direction: "horizontal",
							mouseScrollNavigation:"off",
 							mouseScrollReverse:"default",
							onHoverStop:"on",
							arrows: {
								style:"academia",
								enable:true,
								hide_onmobile:true,
								hide_under:480,
								hide_onleave:false,
								tmp:'',
								left: {
									h_align:"left",
									v_align:"center",
									h_offset:20,
									v_offset:0
								},
								right: {
									h_align:"right",
									v_align:"center",
									h_offset:20,
									v_offset:0
								}
							}
						},
						responsiveLevels:[1240,1024,778,480],
						visibilityLevels:[1240,1024,778,480],
						gridwidth:[1200,1024,778,480],
						gridheight:[700,650,600,600],
						lazyType:"none",
						shadow:0,
						spinner:"spinner0",
						stopLoop:"off",
						stopAfterLoops:-1,
						stopAtSlide:-1,
						shuffle:"off",
						autoHeight:"off",
						disableProgressBar:"on",
						hideThumbsOnMobile:"off",
						hideSliderAtLimit:0,
						hideCaptionAtLimit:0,
						hideAllCaptionAtLilmit:0,
						debugMode:false,
						fallbacks: {
							simplifyAll:"off",
							nextSlideOnWindowFocus:"off",
							disableFocusListener:false,
						}
					});
				}
			});	/*ready*/
		</script>
		<script>
					var htmlDivCss = unescape(".academia.tparrows%20%7B%0A%09cursor%3Apointer%3B%0A%09background%3A%23000%3B%0A%09background%3Argba%280%2C0%2C0%2C0.7%29%3B%0A%09width%3A50px%3B%0A%09height%3A60px%3B%0A%09position%3Aabsolute%3B%0A%09display%3Ablock%3B%0A%09z-index%3A100%3B%0A%20%20%20%20-webkit-transition%3A%20all%20.3s%20%21important%3B%0A%09-moz-transition%3A%20all%20.3s%20%21important%3B%0A%09-o-transition%3A%20all%20.3s%20%21important%3B%0A%09transition%3A%20all%20.3s%20%21important%3B%0A%7D%0A.academia.tparrows%3Ahover%20%7B%0A%09background%3A%23FFBC33%3B%0A%7D%0A.academia.tparrows%3Ahover.tp-leftarrow%3Aafter%0A%7B%0A%09border-top%3A%20solid%2060px%20%23FFBC33%3B%0A%20%20%20%20opacity%3A%201%3B%0A%7D%0A.academia.tparrows%3Ahover.tp-rightarrow%3Aafter%0A%7B%0A%09border-bottom%3A%20solid%2060px%20%23FFBC33%3B%0A%20%20%20%20opacity%3A%201%3B%0A%7D%0A.academia.tparrows%3Abefore%20%7B%0A%09font-family%3A%20%22revicons%22%3B%0A%09font-size%3A18px%3B%0A%20%20%20%20font-weight%3A600%3B%0A%09color%3A%23fff%3B%0A%09display%3Ablock%3B%0A%09line-height%3A%2060px%3B%0A%09text-align%3A%20center%3B%0A%7D%0A.academia.tparrows.tp-leftarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce824%22%3B%0A%7D%0A.academia.tparrows.tp-rightarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce825%22%3B%0A%7D%0A.academia.tparrows%3Aafter%0A%7B%0A%09content%3A%20%27%27%3B%0A%20%20%20%20display%3A%20block%3B%0A%20%20%20%20position%3A%20absolute%3B%0A%20%20%20%20top%3A%200%3B%0A%20%20%20%20bottom%3A%200%3B%0A%20%20%20%20opacity%3A%200.7%3B%0A%20%20%20%20-webkit-transition%3A%20all%20.3s%20%21important%3B%0A%09-moz-transition%3A%20all%20.3s%20%21important%3B%0A%09-o-transition%3A%20all%20.3s%20%21important%3B%0A%09transition%3A%20all%20.3s%20%21important%3B%0A%7D%0A.academia.tparrows.tp-leftarrow%3Aafter%7B%0A%20%20%20%20border-bottom%3A%20solid%200%20transparent%3B%0A%20%20%20%20border-top%3A%20solid%2060px%20%23000000%3B%0A%20%20%20%20border-right%3A%20solid%2010px%20transparent%3B%0A%20%20%20%20left%3A%20100%25%3B%0A%7D%0A.academia.tparrows.tp-rightarrow%3Aafter%7B%0A%09border-bottom%3A%20solid%2060px%20%23000000%3B%0A%20%20%20%20border-top%3A%20solid%200%20transparent%3B%0A%20%20%20%20border-left%3A%20solid%2010px%20transparent%3B%0A%20%20%20%20right%3A%20100%25%3B%0A%7D%0A%0A");
					var htmlDiv = document.getElementById('rs-plugin-settings-inline-css');
					if(htmlDiv) {
						htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
					}
					else{
						var htmlDiv = document.createElement('div');
						htmlDiv.innerHTML = '<style>' + htmlDivCss + '</style>';
						document.getElementsByTagName('head')[0].appendChild(htmlDiv.childNodes[0]);
					}
				  </script>
				</div><!-- END REVOLUTION SLIDER --></div></div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12 vc_hidden-lg vc_hidden-md"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="wpb_revslider_element wpb_content_element">
<div id="rev_slider_6_2_wrapper" class="rev_slider_wrapper fullwidthbanner-container" style="margin:0px auto;background-color:transparent;padding:0px;margin-top:0px;margin-bottom:0px;">
<!-- START REVOLUTION SLIDER 5.2.5 auto mode -->
	<div id="rev_slider_6_2" class="rev_slider fullwidthabanner" style="display:none;" data-version="5.2.5">
<ul>	<!-- SLIDE  -->
	<li data-index="rs-69" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2018/02/Slide-Móvil-100x50.png"  data-delay="8010"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/Slide-Móvil.png"  alt="" title="Slide Móvil"  width="600" height="800" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption rev-btn " 
			 id="slide-69-layer-1" 
			 data-x="['left','left','left','left']" data-hoffset="['177','177','177','177']" 
			 data-y="['top','top','top','top']" data-voffset="['340','340','340','340']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(136, 12, 10, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"https:\/\/www.moralurbanidadycivica.com\/"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			
			style="z-index: 5; white-space: nowrap; font-size: 25px; line-height: 17px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:Roboto;background-color:rgba(0, 0, 0, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);border-radius:3px 3px 3px 3px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">AQUÍ </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-54" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2018/01/movilgraduacion-100x50.jpg"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2018/01/movilgraduacion.jpg"  alt="" title="movilgraduacion"  width="480" height="600" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-54-layer-1" 
			 data-x="['center','center','center','center']" data-hoffset="['1','1','1','103']" 
			 data-y="['top','top','top','top']" data-voffset="['270','270','270','194']" 
						data-width="257"
			data-height="115"
			data-whitespace="normal"
			data-transform_idle="o:1;"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			
			style="z-index: 5; min-width: 257px; max-width: 257px; max-width: 115px; max-width: 115px; white-space: normal; font-size: 45px; line-height: 50px; color: rgba(244, 244, 244, 1.00);text-align:center;">Información Graduación LX </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption rev-btn rev-withicon " 
			 id="slide-54-layer-2" 
			 data-x="['left','left','left','left']" data-hoffset="['172','172','172','291']" 
			 data-y="['top','top','top','top']" data-voffset="['391','391','391','305']" 
						data-width="143"
			data-height="76"
			data-whitespace="normal"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":" http:\/\/www.catolica.edu.sv\/?tribe_events=informacion-graduacion-lx"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			
			style="z-index: 6; min-width: 143px; max-width: 143px; max-width: 76px; max-width: 76px; white-space: normal; font-size: 25px; line-height: 17px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:oswald;background-color:rgba(136, 12, 10, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);border-radius:30px 30px 30px 30px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">Aquí<i class="fa-icon-chevron-right"></i> </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-23" data-transition="curtain-2,boxslide,slidedown" data-slotamount="default,default,default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default,default,default" data-easeout="default,default,default" data-masterspeed="default,default,default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/07/cel-web1-100x50.png"  data-delay="8050"  data-rotate="0,0,0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/07/cel-web1.png"  alt="" title="cel-web1"  width="400" height="680" data-bgposition="center bottom" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-sub-heading-top   tp-resizeme" 
			 id="slide-23-layer-2" 
			 data-x="['left','center','center','center']" data-hoffset="['652','84','-30','-117']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-252','-264','-265','-273']" 
						data-fontsize="['30','28','28','28']"
			data-color="['rgba(66, 66, 66, 1.00)','rgba(0, 21, 255, 1.00)','rgba(0, 21, 255, 1.00)','rgba(49, 52, 73, 1.00)']"
			data-width="['262','none','none','none']"
			data-height="['65','none','none','none']"
			data-whitespace="['normal','nowrap','nowrap','nowrap']"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="649.6875" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.6875" 

			style="z-index: 5; min-width: 262px; max-width: 262px; max-width: 65px; max-width: 65px; white-space: normal; font-size: 30px; color: rgba(66, 66, 66, 1.00);">CONOCE NUESTRO </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-23-layer-1" 
			 data-x="['left','center','center','center']" data-hoffset="['651','232','81','27']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-229','-222','-228','-228']" 
						data-fontsize="['50','60','50','45']"
			data-lineheight="['72','72','72','54']"
			data-color="['rgba(66, 66, 66, 1.00)','rgba(0, 21, 255, 1.00)','rgba(0, 21, 255, 1.00)','rgba(49, 52, 73, 1.00)']"
			data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="899.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 6; white-space: nowrap; font-size: 50px; color: rgba(66, 66, 66, 1.00);">CAMPUS UNICAES </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption academia-sub-heading-bottom   tp-resizeme" 
			 id="slide-23-layer-3" 
			 data-x="['left','center','center','center']" data-hoffset="['714','281','217','76']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-191','-183','-192','-190']" 
						data-color="['rgba(6, 2, 10, 1.00)','rgba(13, 0, 33, 1.00)','rgba(13, 0, 33, 1.00)','rgba(13, 0, 33, 1.00)']"
			data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="x:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;s:1500;e:Power3.easeInOut;" 
			 data-transform_out="y:[100%];s:1010;e:Power4.easeInOut;" 
			 data-mask_in="x:0px;y:0px;s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="1149.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 7; white-space: nowrap; color: rgba(6, 2, 10, 1.00);font-family:Oswald;">Y NUESTRAS CARRERAS UNIVERSITARIAS </div>

		<!-- LAYER NR. 4 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-23-layer-6" 
			 data-x="['left','center','center','center']" data-hoffset="['670','198','142','-96']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-131','-144','-158','-122']" 
						data-fontsize="['16','16','16','25']"
			data-lineheight="['30','22','22','22']"
			data-fontweight="['300','400','400','400']"
			data-color="['rgba(28, 28, 28, 1.00)','rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)']"
			data-width="['141','none','none','none']"
			data-height="none"
			data-whitespace="['normal','nowrap','nowrap','nowrap']"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(255, 255, 255, 1.00);bg:rgba(136, 12, 10, 1.00);"
 
			 data-transform_in="opacity:0;s:1500;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1010;e:Power2.easeInOut;" 
			data-start="1149.84375" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=1057"}]'
			data-responsive_offset="on" 

			 data-end="6989.84375" 

			style="z-index: 8; min-width: 141px; max-width: 141px; white-space: normal; font-size: 16px; line-height: 30px; font-weight: 300; color: rgba(28, 28, 28, 1.00);font-family:Oswald;text-align:center;background-color:rgba(237, 189, 63, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">PREGRADOS </div>

		<!-- LAYER NR. 5 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-23-layer-8" 
			 data-x="['left','center','center','center']" data-hoffset="['835','198','142','120']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-129','-144','-158','-114']" 
						data-fontsize="['16','16','16','25']"
			data-lineheight="['30','22','22','22']"
			data-fontweight="['300','400','400','400']"
			data-color="['rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)','rgba(255, 255, 255, 1.00)','rgba(10, 2, 2, 1.00)']"
			data-width="['141','none','none','177']"
			data-height="['none','none','none','58']"
			data-whitespace="['normal','nowrap','nowrap','normal']"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(10, 0, 2, 1.00);bg:rgba(237, 189, 63, 1.00);"
 
			 data-transform_in="opacity:0;s:1500;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1010;e:Power2.easeInOut;" 
			data-start="1399.6875" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=671"}]'
			data-responsive_offset="on" 

			 data-end="6989.6875" 

			style="z-index: 9; min-width: 141px; max-width: 141px; white-space: normal; font-size: 16px; line-height: 30px; font-weight: 300;font-family:Oswald;text-align:center;background-color:rgba(136, 12, 10, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">POSTGRADOS </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-28" data-transition="slidedown" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/07/cel-web2-100x50.png"  data-delay="7990"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/07/cel-web2.png"  alt="" title="cel-web2"  width="400" height="680" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-28-layer-2" 
			 data-x="['left','left','left','left']" data-hoffset="['84','84','84','84']" 
			 data-y="['top','top','top','top']" data-voffset="['74','74','74','74']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="7590" 

			style="z-index: 5; white-space: nowrap; color: rgba(7, 7, 7, 1.00);">ENTÉRATE DE: </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption rev-btn " 
			 id="slide-28-layer-3" 
			 data-x="['left','left','left','left']" data-hoffset="['157','157','157','146']" 
			 data-y="['top','top','top','top']" data-voffset="['161','161','161','163']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="490" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?post_type=tribe_events"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			 data-end="7620" 

			style="z-index: 6; white-space: nowrap; font-size: 30px; line-height: 17px; font-weight: 500; color: rgba(15, 15, 15, 1.00);font-family:OSWALD;background-color:rgba(237, 189, 63, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">EVENTOS </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption rev-btn " 
			 id="slide-28-layer-4" 
			 data-x="['left','left','left','left']" data-hoffset="['155','155','155','144']" 
			 data-y="['top','top','top','top']" data-voffset="['221','221','221','224']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=861"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			 data-end="7560" 

			style="z-index: 7; white-space: nowrap; font-size: 30px; line-height: 17px; font-weight: 500; color: rgba(255, 255, 255, 1.00);font-family:OSWALD;background-color:rgba(136, 12, 10, 0.75);padding:12px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;cursor:pointer;">NOTICIAS </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-22" data-transition="curtain-1,boxfade,slidedown" data-slotamount="default,default,default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default,default,default" data-easeout="default,default,default" data-masterspeed="default,default,default"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2016/07/unnamed-100x50.jpg"  data-delay="9000"  data-rotate="0,0,0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2016/07/unnamed.jpg"  alt="" title="unnamed"  width="1173" height="782" data-bgposition="right center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption academia-heading   tp-resizeme" 
			 id="slide-22-layer-1" 
			 data-x="['left','left','left','left']" data-hoffset="['71','64','47','27']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-171','-186','-186','-186']" 
						data-fontsize="['60','60','50','30']"
			data-lineheight="['72','72','72','60']"
			data-width="['843','844','844','399']"
			data-height="['145','none','none','none']"
			data-whitespace="normal"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1000;e:Power2.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="700" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="8020" 

			style="z-index: 5; min-width: 843px; max-width: 843px; max-width: 145px; max-width: 145px; white-space: normal; color: rgba(10, 10, 10, 1.00);">CENTRO REGIONAL DE ILOBASCO </div>

		<!-- LAYER NR. 2 -->
		<div class="tp-caption academia-sub-heading   tp-resizeme" 
			 id="slide-22-layer-2" 
			 data-x="['left','left','left','left']" data-hoffset="['72','63','46','29']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-260','-236','-229','-219']" 
						data-fontsize="['65','75','75','35']"
			data-width="['345','339','339','240']"
			data-height="['58','83','83','54']"
			data-whitespace="normal"
			data-transform_idle="o:1;"
 
			 data-transform_in="y:[100%];z:0;rX:0deg;rY:0;rZ:0;sX:1;sY:1;skX:0;skY:0;opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="y:[100%];s:1000;e:Power2.easeInOut;" 
			 data-mask_in="x:0px;y:[100%];s:inherit;e:inherit;" 
			 data-mask_out="x:inherit;y:inherit;s:inherit;e:inherit;" 
			data-start="900" 
			data-splitin="none" 
			data-splitout="none" 
			data-responsive_offset="on" 

			 data-end="8009.8965454102" 

			style="z-index: 6; min-width: 345px; max-width: 345px; max-width: 58px; max-width: 58px; white-space: normal; font-size: 65px; line-height: 50px; color: rgba(10, 10, 10, 1.00);">UNICAES </div>

		<!-- LAYER NR. 3 -->
		<div class="tp-caption academia-button-bg rev-btn  tp-resizeme" 
			 id="slide-22-layer-4" 
			 data-x="['left','left','left','left']" data-hoffset="['399','335','286','215']" 
			 data-y="['middle','middle','middle','middle']" data-voffset="['-140','-125','-129','-116']" 
						data-width="['none','none','none','194']"
			data-height="['none','none','none','77']"
			data-whitespace="['nowrap','nowrap','nowrap','normal']"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(10, 2, 4, 1.00);bg:rgba(237, 189, 63, 1.00);"
 
			 data-transform_in="opacity:0;s:2000;e:Power4.easeInOut;" 
			 data-transform_out="opacity:0;s:1000;e:Power2.easeIn;" 
			data-start="1400" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.cri.catolica.edu.sv\/"}]'
			data-responsive_offset="on" 

			 data-end="7000" 

			style="z-index: 7; white-space: nowrap; font-size: 20px;font-family:Oswald;background-color:rgba(136, 12, 10, 1.00);outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;">Ir al sitio web </div>
	</li>
	<!-- SLIDE  -->
	<li data-index="rs-48" data-transition="fade" data-slotamount="default" data-hideafterloop="0" data-hideslideonmobile="off"  data-easein="default" data-easeout="default" data-masterspeed="300"  data-thumb="http://www.catolica.edu.sv/wp-content/uploads/2017/05/slider-movil-100x50.jpg"  data-delay="7000"  data-rotate="0"  data-saveperformance="off"  data-title="Slide" data-param1="" data-param2="" data-param3="" data-param4="" data-param5="" data-param6="" data-param7="" data-param8="" data-param9="" data-param10="" data-description="">
		<!-- MAIN IMAGE -->
		<img src="http://www.catolica.edu.sv/wp-content/uploads/2017/05/slider-movil.jpg"  alt="" title="slider-movil"  width="480" height="600" data-bgposition="center center" data-bgfit="cover" data-bgrepeat="no-repeat" class="rev-slidebg" data-no-retina>
		<!-- LAYERS -->

		<!-- LAYER NR. 1 -->
		<div class="tp-caption rev-btn rev-hiddenicon " 
			 id="slide-48-layer-1" 
			 data-x="['center','center','center','center']" data-hoffset="['0','0','0','0']" 
			 data-y="['top','top','top','top']" data-voffset="['100','100','100','100']" 
						data-width="none"
			data-height="none"
			data-whitespace="nowrap"
			data-transform_idle="o:1;"
				data-transform_hover="o:1;rX:0;rY:0;rZ:0;z:0;s:0;e:Linear.easeNone;"
				data-style_hover="c:rgba(0, 0, 0, 1.00);bg:rgba(255, 255, 255, 1.00);"
 
			 data-transform_in="opacity:0;s:300;e:Power2.easeInOut;" 
			 data-transform_out="opacity:0;s:300;" 
			data-start="500" 
			data-splitin="none" 
			data-splitout="none" 
			data-actions='[{"event":"click","action":"simplelink","target":"_self","url":"http:\/\/www.catolica.edu.sv\/?page_id=7577"}]'
			data-responsive_offset="on" 
			data-responsive="off"
			
			style="z-index: 5; white-space: nowrap; font-size: 55px; line-height: 20px; font-weight: 900; color: rgba(214, 240, 47, 1.00);font-family:oswald;text-align:center;text-transform:uppercase;background-color:rgba(1, 15, 90, 1.00);padding:25px 35px 12px 35px;border-color:rgba(0, 0, 0, 1.00);border-radius:30px 30px 30px 30px;outline:none;box-shadow:none;box-sizing:border-box;-moz-box-sizing:border-box;-webkit-box-sizing:border-box;letter-spacing:1px;cursor:pointer;">Haz clic <i class="fa-icon-mouse-pointer"></i> </div>
	</li>
</ul>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss="";
						if(htmlDiv) {
							htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
						}else{
							var htmlDiv = document.createElement("div");
							htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
							document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
						}
					</script>
<div class="tp-bannertimer tp-bottom" style="visibility: hidden !important;"></div>	</div>
<script>var htmlDiv = document.getElementById("rs-plugin-settings-inline-css"); var htmlDivCss=".tp-caption.academia-sub-heading-top,.academia-sub-heading-top{color:rgba(255,255,255,1.00);font-size:28px;line-height:33.6px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left}.tp-caption.academia-heading,.academia-heading{color:rgba(255,255,255,1.00);font-size:60px;line-height:72px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left;letter-spacing:0.02em}.tp-caption.academia-sub-heading-bottom,.academia-sub-heading-bottom{color:rgba(255,255,255,1.00);font-size:16px;line-height:19.2px;font-weight:400;font-style:normal;font-family:Roboto;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left}.tp-caption.academia-button-bg,.academia-button-bg{color:rgba(255,255,255,1.00);font-size:12px;line-height:22px;font-weight:400;font-style:normal;font-family:Roboto;padding:11px 30px 11px 30px;text-decoration:none;background-color:rgba(47,167,203,1.00);border-color:transparent;border-style:solid;border-width:0px;border-radius:0px 0px 0px 0px;text-align:left;letter-spacing:0.05em !important;-webkit-transition:all .3s !important;-moz-transition:all .3s !important;-o-transition:all .3s !important;transition:all .3s !important}.tp-caption.academia-button-bg:hover,.academia-button-bg:hover{color:rgba(255,255,255,1.00);text-decoration:none;background-color:rgba(145,95,169,1.00);border-color:transparent;border-style:none;border-width:0px;border-radius:0px 0px 0px 0px}.tp-caption.academia-sub-heading,.academia-sub-heading{color:rgba(255,255,255,1.00);font-size:24px;line-height:28.8px;font-weight:400;font-style:normal;font-family:Oswald;padding:0 0 0 0px;text-decoration:none;background-color:transparent;border-color:transparent;border-style:none;border-width:0px;border-radius:0 0 0 0px;text-align:left;letter-spacing:0.1em}";
				if(htmlDiv) {
					htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
				}else{
					var htmlDiv = document.createElement("div");
					htmlDiv.innerHTML = "<style>" + htmlDivCss + "</style>";
					document.getElementsByTagName("head")[0].appendChild(htmlDiv.childNodes[0]);
				}
			</script>
		<script type="text/javascript">
						/******************************************
				-	PREPARE PLACEHOLDER FOR SLIDER	-
			******************************************/

			var setREVStartSize=function(){
				try{var e=new Object,i=jQuery(window).width(),t=9999,r=0,n=0,l=0,f=0,s=0,h=0;
					e.c = jQuery('#rev_slider_6_2');
					e.responsiveLevels = [1240,1024,778,480];
					e.gridwidth = [1200,1024,778,480];
					e.gridheight = [700,650,600,600];
							
					e.sliderLayout = "auto";
					if(e.responsiveLevels&&(jQuery.each(e.responsiveLevels,function(e,f){f>i&&(t=r=f,l=e),i>f&&f>r&&(r=f,n=e)}),t>r&&(l=n)),f=e.gridheight[l]||e.gridheight[0]||e.gridheight,s=e.gridwidth[l]||e.gridwidth[0]||e.gridwidth,h=i/s,h=h>1?1:h,f=Math.round(h*f),"fullscreen"==e.sliderLayout){var u=(e.c.width(),jQuery(window).height());if(void 0!=e.fullScreenOffsetContainer){var c=e.fullScreenOffsetContainer.split(",");if (c) jQuery.each(c,function(e,i){u=jQuery(i).length>0?u-jQuery(i).outerHeight(!0):u}),e.fullScreenOffset.split("%").length>1&&void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0?u-=jQuery(window).height()*parseInt(e.fullScreenOffset,0)/100:void 0!=e.fullScreenOffset&&e.fullScreenOffset.length>0&&(u-=parseInt(e.fullScreenOffset,0))}f=u}else void 0!=e.minHeight&&f<e.minHeight&&(f=e.minHeight);e.c.closest(".rev_slider_wrapper").css({height:f})
					
				}catch(d){console.log("Failure at Presize of Slider:"+d)}
			};
			
			setREVStartSize();
			
						var tpj=jQuery;
			
			var revapi6;
			tpj(document).ready(function() {
				if(tpj("#rev_slider_6_2").revolution == undefined){
					revslider_showDoubleJqueryError("#rev_slider_6_2");
				}else{
					revapi6 = tpj("#rev_slider_6_2").show().revolution({
						sliderType:"standard",
jsFileLocation:"//www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/js/",
						sliderLayout:"auto",
						dottedOverlay:"none",
						delay:4000,
						navigation: {
							keyboardNavigation:"off",
							keyboard_direction: "horizontal",
							mouseScrollNavigation:"off",
 							mouseScrollReverse:"default",
							onHoverStop:"off",
							arrows: {
								style:"academia",
								enable:true,
								hide_onmobile:true,
								hide_under:480,
								hide_onleave:true,
								hide_delay:200,
								hide_delay_mobile:1200,
								tmp:'',
								left: {
									h_align:"left",
									v_align:"center",
									h_offset:20,
									v_offset:0
								},
								right: {
									h_align:"right",
									v_align:"center",
									h_offset:20,
									v_offset:0
								}
							}
						},
						responsiveLevels:[1240,1024,778,480],
						visibilityLevels:[1240,1024,778,480],
						gridwidth:[1200,1024,778,480],
						gridheight:[700,650,600,600],
						lazyType:"none",
						shadow:0,
						spinner:"spinner0",
						stopLoop:"off",
						stopAfterLoops:-1,
						stopAtSlide:-1,
						shuffle:"off",
						autoHeight:"off",
						disableProgressBar:"on",
						hideThumbsOnMobile:"off",
						hideSliderAtLimit:0,
						hideCaptionAtLimit:0,
						hideAllCaptionAtLilmit:0,
						debugMode:false,
						fallbacks: {
							simplifyAll:"off",
							nextSlideOnWindowFocus:"off",
							disableFocusListener:false,
						}
					});
				}
			});	/*ready*/
		</script>
		<script>
					var htmlDivCss = unescape(".academia.tparrows%20%7B%0A%09cursor%3Apointer%3B%0A%09background%3A%23000%3B%0A%09background%3Argba%280%2C0%2C0%2C0.7%29%3B%0A%09width%3A50px%3B%0A%09height%3A60px%3B%0A%09position%3Aabsolute%3B%0A%09display%3Ablock%3B%0A%09z-index%3A100%3B%0A%20%20%20%20-webkit-transition%3A%20all%20.3s%20%21important%3B%0A%09-moz-transition%3A%20all%20.3s%20%21important%3B%0A%09-o-transition%3A%20all%20.3s%20%21important%3B%0A%09transition%3A%20all%20.3s%20%21important%3B%0A%7D%0A.academia.tparrows%3Ahover%20%7B%0A%09background%3A%23FFBC33%3B%0A%7D%0A.academia.tparrows%3Ahover.tp-leftarrow%3Aafter%0A%7B%0A%09border-top%3A%20solid%2060px%20%23FFBC33%3B%0A%20%20%20%20opacity%3A%201%3B%0A%7D%0A.academia.tparrows%3Ahover.tp-rightarrow%3Aafter%0A%7B%0A%09border-bottom%3A%20solid%2060px%20%23FFBC33%3B%0A%20%20%20%20opacity%3A%201%3B%0A%7D%0A.academia.tparrows%3Abefore%20%7B%0A%09font-family%3A%20%22revicons%22%3B%0A%09font-size%3A18px%3B%0A%20%20%20%20font-weight%3A600%3B%0A%09color%3A%23fff%3B%0A%09display%3Ablock%3B%0A%09line-height%3A%2060px%3B%0A%09text-align%3A%20center%3B%0A%7D%0A.academia.tparrows.tp-leftarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce824%22%3B%0A%7D%0A.academia.tparrows.tp-rightarrow%3Abefore%20%7B%0A%09content%3A%20%22%5Ce825%22%3B%0A%7D%0A.academia.tparrows%3Aafter%0A%7B%0A%09content%3A%20%27%27%3B%0A%20%20%20%20display%3A%20block%3B%0A%20%20%20%20position%3A%20absolute%3B%0A%20%20%20%20top%3A%200%3B%0A%20%20%20%20bottom%3A%200%3B%0A%20%20%20%20opacity%3A%200.7%3B%0A%20%20%20%20-webkit-transition%3A%20all%20.3s%20%21important%3B%0A%09-moz-transition%3A%20all%20.3s%20%21important%3B%0A%09-o-transition%3A%20all%20.3s%20%21important%3B%0A%09transition%3A%20all%20.3s%20%21important%3B%0A%7D%0A.academia.tparrows.tp-leftarrow%3Aafter%7B%0A%20%20%20%20border-bottom%3A%20solid%200%20transparent%3B%0A%20%20%20%20border-top%3A%20solid%2060px%20%23000000%3B%0A%20%20%20%20border-right%3A%20solid%2010px%20transparent%3B%0A%20%20%20%20left%3A%20100%25%3B%0A%7D%0A.academia.tparrows.tp-rightarrow%3Aafter%7B%0A%09border-bottom%3A%20solid%2060px%20%23000000%3B%0A%20%20%20%20border-top%3A%20solid%200%20transparent%3B%0A%20%20%20%20border-left%3A%20solid%2010px%20transparent%3B%0A%20%20%20%20right%3A%20100%25%3B%0A%7D%0A%0A");
					var htmlDiv = document.getElementById('rs-plugin-settings-inline-css');
					if(htmlDiv) {
						htmlDiv.innerHTML = htmlDiv.innerHTML + htmlDivCss;
					}
					else{
						var htmlDiv = document.createElement('div');
						htmlDiv.innerHTML = '<style>' + htmlDivCss + '</style>';
						document.getElementsByTagName('head')[0].appendChild(htmlDiv.childNodes[0]);
					}
				  </script>
				</div><!-- END REVOLUTION SLIDER --></div></div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12 vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center mg-top-100 mg-bottom-60" >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    MENSAJE DEL RECTOR                </h2>
                                <p class="fs-14">
                    BIENVENIDOS                </p>
                            </div>
            </div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-4 vc_hidden-lg vc_hidden-md"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<div class="heading color-dark text-center mg-bottom-60">
<p><img class="alignnone size-full wp-image-4185" src="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" alt="estrellas" width="56" height="25" /></p>
<h2 class="heading-color fs-38">UNIVERSIDAD CATÓLICA DE EL SALVADOR</h2>
</div>

		</div>
	</div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h3 style="text-align: center;">BIENVENIDOS</h3>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<hr />
<h4 style="text-align: center;"><strong>Mensaje del rector</strong></h4>
<hr />

		</div>
	</div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<div class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Rector-8x12-web-321x482.jpg" width="321" height="482" alt="Rector-8x12-web" title="Rector-8x12-web" /></div>
		</figure>
	</div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: justify;">Hay dos tareas esenciales para cualquier universidad: la primera, consiste en conseguir una educación profesional óptima para los alumnos, adquirir un prestigio institucional en términos de capacitación profesional y formación; la otra tarea, más difícil, es la formación del ser humano.<br />
Si repasamos la historia vemos cómo las universidades eran realmente elementos de formación de la cultura europea. Ahora tenemos otra vez la misma oportunidad, máxime dentro del modelo competitivo que internacionalmente se ha impuesto. Para ser el mejor, cada uno en su campo, ha de estar en continua comunicación y cooperación con otras universidades del resto del mundo. Esta internacionalización es una gran oportunidad, algo muy bueno.<br />
Al mismo tiempo, la formación integral del ser humano, aspecto crucial, va en camino de perderse, a no ser que alguno de aquellos que conocen su importancia busquen cómo fomentarla de nuevo. Y eso sólo puede hacerse partiendo de la premisa básica de que la universidad no es un negocio como cualquier otro.</p>

		</div>
	</div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: justify;">De algún modo, nosotros tenemos que enseñar a la sociedad un modelo nuevo. Debemos decir: &#8220;esta es la identidad de la universidad&#8221;. Nosotros formamos al ser humano, además de darle una educación estrictamente profesional: es la buena conjunción de estos dos factores la que es capaz de hacer feliz al hombre. Debemos saber quiénes somos, la trascendental tarea que estamos llamados a cumplir, y esto lo descubriremos sólo si, olvidándonos momentáneamente del modelo utilitarista, nos paramos a leer un poco de filosofía y ética.</p>
<p style="text-align: justify;">Las ansias de saber lo que uno es son, paradójicamente, mucho mayores hoy que en otros momentos históricos, a pesar de que nuestras condiciones materiales de vida desbordan con mucho aquellas que nuestros antecesores podían soñar.</p>
<p>&nbsp;</p>
<p style="text-align: right;">Mons. Miguel Ángel Morán Aquino<br />
Palabras en la LIX Graduación UNICAES</p>

		</div>
	</div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid vc_custom_1518622494109"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="https://www.moralurbanidadycivica.com/" target="_blank" class="vc_single_image-wrapper   vc_box_border_grey"><img width="1317" height="310" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_Sitio_UNICAES.png" class="vc_single_image-img attachment-full" alt="" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_Sitio_UNICAES.png 1317w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_Sitio_UNICAES-300x71.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_Sitio_UNICAES-1024x241.png 1024w" sizes="(max-width: 1317px) 100vw, 1317px" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div>
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<div class="heading color-dark text-center mg-bottom-60">
<p><img class="alignnone size-full wp-image-4185" src="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" alt="estrellas" width="56" height="25" /></p>
<h2 class="heading-color fs-38"><a style="color: #000000;" href="http://www.catolica.edu.sv/?page_id=7577">ENTÉRATE DE LOS PROCESOS</a></h2>
</div>

		</div>
	</div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://www.catolica.edu.sv/?page_id=7577" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img width="1024" height="512" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/UNICAES-EN-LINEA-BOTON-1024x512.jpg" class="vc_single_image-img attachment-large" alt="" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/UNICAES-EN-LINEA-BOTON-1024x512.jpg 1024w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/UNICAES-EN-LINEA-BOTON-300x150.jpg 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/UNICAES-EN-LINEA-BOTON.jpg 1200w" sizes="(max-width: 1024px) 100vw, 1024px" /></a>
		</figure>
	</div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-6"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center mg-top-100 mg-bottom-60" >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Facultad Multidisciplinaria                </h2>
                                <p class="fs-14">
                     de Ilobasco                </p>
                            </div>
            <div class="vc_btn3-container vc_btn3-center"><a class="vc_general vc_btn3 vc_btn3-size-lg vc_btn3-shape-rounded vc_btn3-style-3d vc_btn3-block vc_btn3-icon-left vc_btn3-color-peacoc" href="http://www.cri.catolica.edu.sv" title="FACULTAD MULTIDISCIPLINARIA DE ILOBASCO" target="_blank"><i class="vc_btn3-icon fa fa-home"></i> Ir al sitio UNICAES Ilobasco</a></div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-6"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center mg-top-100 mg-bottom-60" >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Servicios Académicos                </h2>
                                <p class="fs-14">
                     Registro Académico                </p>
                            </div>
            <div class="vc_btn3-container vc_btn3-center"><a class="vc_general vc_btn3 vc_btn3-size-lg vc_btn3-shape-rounded vc_btn3-style-3d vc_btn3-block vc_btn3-icon-left vc_btn3-color-primary" href="http://www.registroacademico.catolica.edu.sv" title="Registro Académico UNICAES" target="_blank"><i class="vc_btn3-icon fa fa-home"></i> Ir al sitio Registro Académico</a></div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center mg-top-100 mg-bottom-60" >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Servicios Online                </h2>
                            </div>
            </div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 30px" ><span class="vc_empty_space_inner"></span></div>
<div class="wpb_gallery wpb_content_element vc_clearfix"><div class="wpb_wrapper"><div class="wpb_gallery_slides wpb_flexslider flexslider_fade flexslider" data-interval="3" data-flex_fx="fade"><ul class="slides"><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/photo-web4.png" width="800" height="600" alt="photo-web4" title="photo-web4" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/photo-web5.png" width="800" height="600" alt="photo-web5" title="photo-web5" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/photo-web1.png" width="800" height="600" alt="photo-web1" title="photo-web1" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/photo-web7.png" width="800" height="600" alt="photo-web7" title="photo-web7" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/photo-web6.png" width="800" height="600" alt="photo-web6" title="photo-web6" /></li></ul></div></div></div></div></div></div><div class="wpb_column vc_column_container vc_col-sm-6"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 32px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-3"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://www.catolica.edu.sv/?page_id=2935" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/moodle-75x75.jpg" width="75" height="75" alt="moodle UNICAES" title="moodle UNICAES" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://mail.google.com/a/catolica.edu.sv/" target="_blank" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/mail-1-75x75.png" width="75" height="75" alt="Email" title="Email" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://www.catalogo.catolica.edu.sv" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/catalogoth2014-75x75.jpg" width="75" height="75" alt="Biblioteca" title="Biblioteca" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://search.ebscohost.com/Community.aspx?authtype=ip&amp;ugt=723731463C9635073786355632853E7228E368D36813669366E320E330133603&amp;IsAdminMobile=N&amp;encid=22D731163C5635373736357632353C47385378C378C376C376C370C370C376C33013" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/EBSCO-75x75.png" width="75" height="75" alt="EBSCO" title="EBSCO" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-9"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=2935"><span style="color: #800000;">AULAS VIRTUALES</span></a></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: center;"><a href="http://www.moodle.catolica.edu.sv/moodle/" target="_blank" rel="noopener noreferrer">Presenciales</a> &#8211; <a href="http://www.moodle.catolica.edu.sv/moodlesp/" target="_blank" rel="noopener noreferrer">Semi-presenciales</a> &#8211; <a href="http://www.catolica.edu.sv/?page_id=4236" target="_blank" rel="noopener noreferrer">Postgrados</a></p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 25px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://mail.google.com/a/catolica.edu.sv/" target="_blank" rel="noopener noreferrer">CORREO ELECTRÓNICO</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: center;"><a href="https://www.sistemas2.catolica.edu.sv" class="broken_link">Crea tu correo institucional</a><br />
<a href="http://mail.google.com/a/catolica.edu.sv/">Ingresa a tu correo institucional</a> (@catolica.edu.sv)</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 20px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://www.catalogo.catolica.edu.sv">CATÁLOGO EN LÍNEA</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: center;">Consulta y reserva de libros de Biblioteca Miguel de Cervantes.</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 25px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://search.ebscohost.com/Community.aspx?authtype=ip&amp;ugt=723731463C9635073786355632853E7224E368D36813669366E320E330133603&amp;IsAdminMobile=N&amp;encid=22D731263C3635973756359632953C97349378C378C376C376C370C370C376C33013&amp;selectServicesToken=AxkK4bDrwP6YERmOqJeg-pJBQm-Z8-ZXj0etBvg1v5_0F0PlRd0mQfb6bt_OgeNJE19EQfMrIRM5S3TpETz7uO3DcsbM0fbSQXZHZs1hOY_t_pKBObvi-SgbxOUnf9zVZbVjXqaLecQDheK_wiQh1zace1vGX3SDIoJBRdcCdke7ZKF10iAuKNpjeaG8rLGT5zuPiw8dysHtHrZpIGLAg0TCRznlPe7aOn-U4OHSZDAr-jGxKXfs9cckUvlhh_qpZxMtsrXpAZZks9wZ8Nf3UxSDKA">EBSCO</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: center;">EBSCO es una base de datos que ofrece textos completos, índices y publicaciones periódicas académicas</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 20px" ><span class="vc_empty_space_inner"></span></div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div></div></div></div><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper"></div></div></div></div></div><div class="vc_empty_space"  style="height: 72px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-lg vc_hidden-md vc_hidden-sm vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="wpb_gallery wpb_content_element vc_clearfix"><div class="wpb_wrapper"><div class="wpb_gallery_slides wpb_flexslider flexslider_fade flexslider" data-interval="3" data-flex_fx="fade"><ul class="slides"><li></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/IMG_0175-compressor-1000x700.jpg" width="1000" height="700" alt="IMG_0175-compressor" title="IMG_0175-compressor" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/pag.95-anuario-1024x683-compressor-1000x700.jpg" width="1000" height="700" alt="pag.95-anuario-1024x683-compressor" title="pag.95-anuario-1024x683-compressor" /></li><li><img class="" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/IMG_9539-compressor-1000x700.jpg" width="1000" height="700" alt="IMG_9539-compressor" title="IMG_9539-compressor" /></li></ul></div></div></div></div></div></div><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-lg vc_hidden-md vc_hidden-sm vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-3"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://172.18.0.219/?page_id=2935" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/moodle-75x75.jpg" width="75" height="75" alt="moodle UNICAES" title="moodle UNICAES" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://search.ebscohost.com/Community.aspx?authtype=ip&amp;ugt=723731463C9635073786355632853E7228E368D36813669366E320E330133603&amp;IsAdminMobile=N&amp;encid=22D731163C5635373736357632353C47385378C378C376C376C370C370C376C33013" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/EBSCO-75x75.png" width="75" height="75" alt="EBSCO" title="EBSCO" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://gmail.com" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/mail-1-75x75.png" width="75" height="75" alt="Email" title="Email" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://www.catalogo.catolica.edu.sv" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/05/catalogoth2014-75x75.jpg" width="75" height="75" alt="Biblioteca" title="Biblioteca" /></a>
		</figure>
	</div>
<div class="vc_empty_space"  style="height: 15px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_single_image wpb_content_element vc_align_center">
		
		<figure class="wpb_wrapper vc_figure">
			<a href="http://172.18.0.219/?page_id=2110" target="_self" class="vc_single_image-wrapper   vc_box_border_grey"><img class="vc_single_image-img " src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Notas-75x75.png" width="75" height="75" alt="Notas" title="Notas" /></a>
		</figure>
	</div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-9"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=2935"><span style="color: #800000;">AULAS VIRTUALES</span></a></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="text-align: center;"><span style="color: #808080;"><span style="text-decoration: underline;"><a style="color: #808080; text-decoration: underline;" href="http://www.moodle.catolica.edu.sv/moodle/" target="_blank" rel="noopener noreferrer">Presenciales</a></span>  <span style="text-decoration: underline;"><a style="color: #808080; text-decoration: underline;" href="http://www.moodle.catolica.edu.sv/moodlesp/" target="_blank" rel="noopener noreferrer">Semi-presenciales</a></span>  <span style="text-decoration: underline;"><a style="color: #808080; text-decoration: underline;" href="http://www.catolica.edu.sv/?page_id=4236" target="_blank" rel="noopener noreferrer">Postgrados</a></span></span></p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 20px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://search.ebscohost.com/Community.aspx?authtype=ip&amp;ugt=723731463C9635073786355632853E7224E368D36813669366E320E330133603&amp;IsAdminMobile=N&amp;encid=22D731263C3635973756359632953C97349378C378C376C376C370C370C376C33013&amp;selectServicesToken=AxkK4bDrwP6YERmOqJeg-pJBQm-Z8-ZXj0etBvg1v5_0F0PlRd0mQfb6bt_OgeNJE19EQfMrIRM5S3TpETz7uO3DcsbM0fbSQXZHZs1hOY_t_pKBObvi-SgbxOUnf9zVZbVjXqaLecQDheK_wiQh1zace1vGX3SDIoJBRdcCdke7ZKF10iAuKNpjeaG8rLGT5zuPiw8dysHtHrZpIGLAg0TCRznlPe7aOn-U4OHSZDAr-jGxKXfs9cckUvlhh_qpZxMtsrXpAZZks9wZ8Nf3UxSDKA">EBSCO</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p>EBSCO es una base de datos que ofrece textos completos, índices y publicaciones periódicas académicas</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 20px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://gmail.com">CORREO ELECTRÓNICO</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p>Correo institucional (@catolica.edu.sv), Drive (almacenamiento ilimitado)</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 20px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://www.catalogo.catolica.edu.sv">CATÁLOGO EN LÍNEA</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 5px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p>Consulta y reserva de libros de Biblioteca Miguel de Cervantes.</p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 30px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h4 style="text-align: center;"><span style="color: #800000;"><a style="color: #800000;" href="http://www.catolica.edu.sv/?page_id=2110">HISTORIAL DE NOTAS</a></span></h4>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div>
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p>Consulta tus notas de cada ciclo académico, crea tu correo institucional y cambia la contraseña inicial.</p>

		</div>
	</div>
</div></div></div></div></div><div class="vc_empty_space"  style="height: 72px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid mg-bottom-40"><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center " >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Calendario Académico                </h2>
                            </div>
            <div class="vc_empty_space"  style="height: 18px" ><span class="vc_empty_space_inner"></span></div>
<div class="vc_btn3-container vc_btn3-center"><a class="vc_general vc_btn3 vc_btn3-size-lg vc_btn3-shape-rounded vc_btn3-style-modern vc_btn3-block vc_btn3-icon-left vc_btn3-color-peacoc" href="http://www.catolica.edu.sv/wp-content/uploads/2017/12/CALENDARIO-ACADÉMICO-2018-version-final-130717.pdf" title="Calendario Academico" target="_blank"><i class="vc_btn3-icon fa fa-calendar"></i> Descárgalo</a></div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center " >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Oportunidades                </h2>
                            </div>
            <div class="vc_empty_space"  style="height: 18px" ><span class="vc_empty_space_inner"></span></div>
<div class="vc_btn3-container vc_btn3-center"><a class="vc_general vc_btn3 vc_btn3-size-lg vc_btn3-shape-rounded vc_btn3-style-modern vc_btn3-block vc_btn3-icon-left vc_btn3-color-blue" href="http://www.catolica.edu.sv/?page_id=5994" title="Oportunidades" target="_blank"><i class="vc_btn3-icon fa fa-book"></i> Entérate</a></div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-4"><div class="vc_column-inner "><div class="wpb_wrapper">            <div class="heading color-dark text-center " >
                                    <span class="s-color"><i class="fa fa-star"></i></span>
                                                <h2 class="heading-color fs-38">
                    Anuario Académico                </h2>
                            </div>
            <div class="vc_empty_space"  style="height: 18px" ><span class="vc_empty_space_inner"></span></div>
<div class="vc_btn3-container vc_btn3-center"><a class="vc_general vc_btn3 vc_btn3-size-lg vc_btn3-shape-rounded vc_btn3-style-modern vc_btn3-block vc_btn3-icon-left vc_btn3-color-primary" href="https://drive.google.com/open?id=1i4LjSK3rXF_0UzsP3qXbLk5r-RPDTxkd" title="Anuario Academico" target="_blank"><i class="vc_btn3-icon fa fa-book"></i> Descárgalo</a></div>
</div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid mg-bottom-40"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<div class="heading color-dark text-center mg-bottom-60">
<p><img class="alignnone size-full wp-image-4185" src="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" alt="estrellas" width="56" height="25" /></p>
<h2 class="heading-color fs-38"><a style="color: #000000;" href="http://www.catolica.edu.sv/?page_id=861">Últimas Noticias</a></h2>
</div>

		</div>
	</div>
            <div class="shortcode-blog-wrap  " >
                <div class="blog-wrap grid">
                    <div class="blog-inner clearfix blog-style-grid no-sidebar blog-col-3">
                        
<article id="post-9568" class="clearfix post-9568 post type-post status-publish format-gallery hentry category-noticias post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2262-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2262-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2287-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2287-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2308-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2308-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2288-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2288-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2275-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2275-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2291-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2291-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2327-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2327-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2339-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2339-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2286-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2286-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2320-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2320-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2344-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2344-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2330-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2330-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9568" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2345-1024x768-570x570.jpg" alt="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9568]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A2345-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9568" rel="bookmark" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017"> 14 marzo, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9568" rel="bookmark" title="Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017">Justicia y transparencia: rendición de cuentas de becas y estipendios MINED 2017</a>
        </h3>
        <div class="entry-excerpt">
            “Un acto de justicia y transparencia”, así calificó el Vicerrector Regional de UNICAES, Monseñor Fray Elías Rauda, a la ceremonia de rendición de cuentas del proyecto "Becas y estipendios MINED para educación técnica superior", administrado por el Centro Regional de Ilobasco, durante el 2017. Al evento asistieron representantes del Ministerio de Educación, autoridades universitarias y [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9568#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    350            </li>
        </ul>        </div>
    </div>
</article>



<article id="post-9536" class="clearfix post-9536 post type-post status-publish format-gallery hentry category-noticias post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9536" title="Noticias UNICAES en La Prensa Gráfica &#8211; Marzo" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/lpg-marzo-2018-570x570.png" alt="Noticias UNICAES en La Prensa Gráfica &#8211; Marzo" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9536]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/lpg-marzo-2018.png" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9536" rel="bookmark" title="Noticias UNICAES en La Prensa Gráfica &#8211; Marzo"> 10 marzo, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9536" rel="bookmark" title="Noticias UNICAES en La Prensa Gráfica &#8211; Marzo">Noticias UNICAES en La Prensa Gráfica &#8211; Marzo</a>
        </h3>
        <div class="entry-excerpt">
            VER PUBLICACIÓN DE MARZO AQUÍ Este mes, en La Prensa Gráfica, publicamos la investigación dulce de la vainilla, donde investigadores del Laboratorio de Tejidos y Cultivos vegetales de UNICAES, nos comparten algunos de sus resultados científicos, así como los beneficios e impacto de este producto agrícola en la economía de El Salvador. También, te contamos [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9536#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    511            </li>
        </ul>        </div>
    </div>
</article>



<article id="post-9517" class="clearfix post-9517 post type-post status-publish format-gallery hentry category-noticias post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A0002-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A0002.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9834-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9834.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9853-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9853.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9897-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9897.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9906-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9906.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9913-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9913.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9923-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9923.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9946-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9946.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9517" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9958-570x570.jpg" alt="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9517]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9958.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9517" rel="bookmark" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR"> 7 marzo, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9517" rel="bookmark" title="ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR">ALEMANIA, UN PAÍS Y UN IDIOMA POR EXPLORAR</a>
        </h3>
        <div class="entry-excerpt">
            En su estadía por UNICAES, el joven investigador de Alemania ha compartido parte de su trabajo de doctorado, con estudiantes de UNICAES. Desde hace dos semanas, en UNICAES nos visita el profesor de literatura española, Tim Christmann, de la Universidad de Saarland, Alemania. El propósito de su estadía es compartir experiencias culturales y científicas de [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9517#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    118            </li>
        </ul>        </div>
    </div>
</article>



<article id="post-9508" class="clearfix post-9508 post type-post status-publish format-gallery hentry category-noticias post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9508" title="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9805-570x570.jpg" alt="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9508]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9805.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9508" title="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9809-570x570.jpg" alt="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9508]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9809.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9508" title="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9828-570x570.jpg" alt="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9508]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/03/0A8A9828.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9508" rel="bookmark" title="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA"> 1 marzo, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9508" rel="bookmark" title="VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA">VAINILLA, UNA INVESTIGACIÓN DULCE PARA EL PALADAR CIENTÍFICO EN AGRONOMÍA</a>
        </h3>
        <div class="entry-excerpt">
            A simple vista, la vainilla es una planta poco atractiva; incluso, hasta puede pasar desapercibida, pero lo que muchos ignoran es que la vainilla es una orquídea única dentro de su género, con gran potencial económico en la industria agronómica y productiva de una nación. O por lo menos, así concluye la investigación “Germinación in vitro [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9508#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    1795            </li>
        </ul>        </div>
    </div>
</article>



<article id="post-9387" class="clearfix post-9387 post type-post status-publish format-gallery hentry category-noticias post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1368-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1368.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A7623-1024x768-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A7623-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1374-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1374.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1365-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1365.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A0678-1024x768-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A0678-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1372-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1372.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1367-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1367.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A0674-1024x768-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/0A8A0674-1024x768.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9387" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1370-570x570.jpg" alt="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9387]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG_1370.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9387" rel="bookmark" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL"> 9 febrero, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9387" rel="bookmark" title="MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL">MAESTRÍAS UNICAES: CASOS DE ÉXITO PROFESIONAL</a>
        </h3>
        <div class="entry-excerpt">
            Una oportunidad de superación profesional es la que se puede tener estudiando una maestría o un programa de especialización académica; UNICAES, como parte de sus prácticas de formación continua y de actualización del conocimiento, facilita cuatro maestrías en diferentes áreas de estudio. Deseo de superación profesional, satisfacción personal o, simplemente, el ímpetu por cultivar y [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9387#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    881            </li>
        </ul>        </div>
    </div>
</article>



<article id="post-9374" class="clearfix post-9374 post type-post status-publish format-gallery hentry category-fac-de-cc-de-salud category-noticias tag-bioseguridad tag-doctorado-en-medicina tag-facultad-ciencias-de-la-salud tag-oms tag-santa-ana post_format-post-format-gallery">
            <div class="entry-thumbnail-wrap">
            <div class='owl-carousel' data-plugin-options='{"items" : 1, "dots" : false, "nav" : true, "animateOut" : "fadeOut", "animateIn" : "fadeIn", "autoplay" : true, "loop" : false}'><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9374" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0002-570x570.jpg" alt="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9374]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0002.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9374" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0003-570x570.jpg" alt="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9374]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0003.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9374" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0005-570x570.jpg" alt="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9374]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0005.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9374" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0006-570x570.jpg" alt="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9374]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0006.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div><div class="entry-thumbnail">
                        <a href="http://www.catolica.edu.sv/?p=9374" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" class="entry-thumbnail-overlay">
                            <img width="570" height="570" class="img-responsive" src="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0007-570x570.jpg" alt="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE" />
                        </a>
                        <a data-rel="prettyPhoto[blog_9374]" href="http://www.catolica.edu.sv/wp-content/uploads/2018/02/IMG-20180205-WA0007.jpg" class="prettyPhoto"><i class="fa fa-expand"></i></a>
                      </div></div>                            <div class="entry-format-date">
                    <span class="entry-icon-format">
                        <i class="fa fa-file-image-o"></i>
                    </span>
                    <span class="entry-date">
                        <a href="http://www.catolica.edu.sv/?p=9374" rel="bookmark" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE"> 8 febrero, 2018 </a>
                    </span>
                </div>
                    </div>
        <div class="entry-content-wrap">
        <h3 class="entry-post-title p-font">
            <a href="http://www.catolica.edu.sv/?p=9374" rel="bookmark" title="CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE">CURSO DE BIOSEGURIDAD: PARA UNA ATENCIÓN MÁS SEGURA DEL PACIENTE</a>
        </h3>
        <div class="entry-excerpt">
            De acuerdo con la Organización Mundial de la Salud (OMS), para garantizar la seguridad del paciente en una intervención clínica o quirúrgica, se deben contemplar algunos pasos esenciales en materia de higiene y limpieza. En esta sintonía, la Facultad de Ciencias de la Salud de UNICAES, organizó el 3° Curso de Bioseguridad, con el objetivo [...]        </div>
        <div class="entry-post-meta-wrap">
            <ul class="entry-meta s-font">
    <li class="entry-meta-author">
        <i class="fa fa-user"></i>
        <a href="http://www.catolica.edu.sv/?author=2">Unidad de Comunicaciones y Mercadeo</a>    </li>

            <li class="entry-meta-comment">
            <a href="http://www.catolica.edu.sv/?p=9374#respond"><i class="fa fa-comments"></i> 0</a>        </li>
        <li class="entry-meta-view">
        <i class="fa fa-eye"></i>
                    460            </li>
        </ul>        </div>
    </div>
</article>


                    </div>

                                            <div class="blog-paging-default">
                            <ul class='pagination'>
	<li><a class="next page-numbers" href="http://www.catolica.edu.sv/?paged=2"><span>Next</span></a></li>
	<li><span class='page-numbers current'>1</span></li>
	<li><a class='page-numbers' href='http://www.catolica.edu.sv/?paged=2'>2</a></li>
	<li><span class="page-numbers dots">&hellip;</span></li>
	<li><a class='page-numbers' href='http://www.catolica.edu.sv/?paged=28'>28</a></li>
</ul>
                        </div>
                    
                </div>
            </div>
            </div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-6"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-9"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><span style="color: #1e73be;">Acreditaciones </span></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div>
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p><img class="aligncenter wp-image-2004" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras-300x269.png" alt="CdA letras negras" width="150" height="134" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras-300x269.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras.png 343w" sizes="(max-width: 150px) 100vw, 150px" /></p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 32px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=3419">Asociaciones y Redes</a></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 12px" ><span class="vc_empty_space_inner"></span></div>
<div class="vc_empty_space"  style="height: 32px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div>
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignnone wp-image-6770 size-full" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices.jpg" alt="" width="144" height="95" /></a><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignnone wp-image-6762 size-full" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cca.jpg" alt="" width="112" height="94" /></a></p>
<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignleft wp-image-6748" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/LOGO-AUPRIDES-v11-300x274.png" alt="" width="104" height="95" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/LOGO-AUPRIDES-v11-300x274.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/LOGO-AUPRIDES-v11.png 398w" sizes="(max-width: 104px) 100vw, 104px" /></a></p>
<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignnone wp-image-6768 size-full" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype1.jpg" alt="" width="107" height="47" /></a></p>
<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="wp-image-6763 size-full alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro.jpg" alt="" width="144" height="96" /></a><img class="alignnone size-medium wp-image-7869" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-ODUCAL-Fondo-Transparente1-300x80.png" alt="" width="300" height="80" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-ODUCAL-Fondo-Transparente1-300x80.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-ODUCAL-Fondo-Transparente1.png 581w" sizes="(max-width: 300px) 100vw, 300px" /></p>
<p style="padding-left: 60px;"><img class="alignnone size-full wp-image-9428" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Catholic-Higher-Education.png" alt="" width="200" height="222" /><img class="alignnone size-medium wp-image-9423" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo-HACU-144x300.gif" alt="" width="144" height="300" /></p>

		</div>
	</div>
</div></div></div><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-md vc_hidden-sm vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=3347">Internacionalización</a></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 12px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="padding-left: 90px;"><img class="size-medium wp-image-8304 alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_UPAEP-300x78.png" alt="" width="300" height="78" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_UPAEP-300x78.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/Logo_UPAEP.png 615w" sizes="(max-width: 300px) 100vw, 300px" /><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="wp-image-3399 alignright" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/AmityInstitute.png" alt="amityinstitute" width="218" height="156" /><img class="size-medium wp-image-8303 alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-vector-universidad-navarra-300x152.jpg" alt="" width="300" height="152" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-vector-universidad-navarra-300x152.jpg 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-vector-universidad-navarra.jpg 630w" sizes="(max-width: 300px) 100vw, 300px" /></a><img class="size-medium wp-image-8305 alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/neiu_wordmark_color-300x51.jpg" alt="" width="300" height="51" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/neiu_wordmark_color-300x51.jpg 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/neiu_wordmark_color-1024x175.jpg 1024w" sizes="(max-width: 300px) 100vw, 300px" /></p>
<p style="text-align: justify; padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="wp-image-8306 size-thumbnail alignnone" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg-150x150.png" alt="" width="150" height="150" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg-150x150.png 150w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg-300x300.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg-1024x1024.png 1024w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/1200px-Logo_Masaryk_University.svg.png 1200w" sizes="(max-width: 150px) 100vw, 150px" /><img class="aligncenter wp-image-3400 size-thumbnail" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-150x150.png" alt="memorialuniversityofnewfoundlandlogo" width="150" height="150" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-150x150.png 150w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-300x300.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo.png 400w" sizes="(max-width: 150px) 100vw, 150px" /></a></p>
<p><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="wp-image-3396 alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-300x61.png" alt="logo-erasmus-plus" width="260" height="53" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-300x61.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-1024x209.png 1024w" sizes="(max-width: 260px) 100vw, 260px" /></a><img class="wp-image-2011 alignright" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-300x74.png" alt="university-of-alberta-logo" width="268" height="66" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-300x74.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-768x190.png 768w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo.png 1000w" sizes="(max-width: 268px) 100vw, 268px" /><br />
<a href="http://www.catolica.edu.sv/?page_id=3347"><img class="wp-image-3397 alignleft" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-300x130.png" alt="uppsalalogo" width="258" height="112" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-300x130.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-1024x443.png 1024w" sizes="(max-width: 258px) 100vw, 258px" /></a><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="wp-image-3398 alignright" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen-300x150.png" alt="coop_externa-rrii_2016-02-26_becas_canada_elap_imagen" width="276" height="138" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen-300x150.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen.png 600w" sizes="(max-width: 276px) 100vw, 276px" /></a></p>

		</div>
	</div>
</div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-lg vc_hidden-md vc_hidden-sm vc_hidden-xs"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="fullwidth" ><div class="vc_row wpb_row vc_inner vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-9"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=3416">Acreditaciones</a></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div>
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="aligncenter wp-image-2004" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras-300x269.png" alt="CdA letras negras" width="150" height="134" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras-300x269.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/CdA-letras-negras.png 343w" sizes="(max-width: 150px) 100vw, 150px" /></a></p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 32px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=3419">Asociaciones y Redes</a></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 12px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignleft wp-image-2006" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices-1-300x248.jpg" alt="raices" width="114" height="94" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices-1-300x248.jpg 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices-1-768x635.jpg 768w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/raices-1.jpg 886w" sizes="(max-width: 114px) 100vw, 114px" /></a><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignnone wp-image-2008" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/ccaa-300x252.png" alt="ccaa" width="112" height="94" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/ccaa-300x252.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/ccaa.png 380w" sizes="(max-width: 112px) 100vw, 112px" /></a></p>
<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3419"><img class="alignleft wp-image-2009" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype-300x264.png" alt="cdmype" width="107" height="94" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype-300x264.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/cdmype.png 362w" sizes="(max-width: 107px) 100vw, 107px" /><img class="alignnone wp-image-2007" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro-300x199.png" alt="innovagro" width="144" height="95" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro-300x199.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/innovagro.png 481w" sizes="(max-width: 144px) 100vw, 144px" /></a></p>

		</div>
	</div>
<div class="vc_empty_space"  style="height: 32px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div></div></div></div><div class="wpb_column vc_column_container vc_col-sm-6 vc_hidden-lg vc_hidden-md"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h1 style="text-align: center;"><a href="http://www.catolica.edu.sv/?page_id=3347">Internacionalización</a></h1>

		</div>
	</div>
<div class="vc_separator wpb_content_element vc_separator_align_center vc_sep_width_100 vc_sep_shadow vc_sep_pos_align_center vc_separator_no_text"><span class="vc_sep_holder vc_sep_holder_l"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span><span class="vc_sep_holder vc_sep_holder_r"><span  style="border-color:#880c0a;" class="vc_sep_line"></span></span>
</div><div class="vc_empty_space"  style="height: 12px" ><span class="vc_empty_space_inner"></span></div>

	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<p><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="alignleft wp-image-3399" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/AmityInstitute.png" alt="amityinstitute" width="218" height="156" /></a></p>
<p style="text-align: justify; padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="alignnone wp-image-3400" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-300x300.png" alt="memorialuniversityofnewfoundlandlogo" width="145" height="145" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-300x300.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo-150x150.png 150w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/MemorialUniversityofNewfoundlandlogo.png 400w" sizes="(max-width: 145px) 100vw, 145px" /></a></p>
<p style="padding-left: 60px;"><a href="http://www.catolica.edu.sv/?page_id=3347"><img class="alignnone wp-image-3396" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-300x61.png" alt="logo-erasmus-plus" width="260" height="53" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-300x61.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/logo-erasmus-plus-1024x209.png 1024w" sizes="(max-width: 260px) 100vw, 260px" /></a><img class="alignnone wp-image-2011" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-300x74.png" alt="university-of-alberta-logo" width="268" height="66" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-300x74.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo-768x190.png 768w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/university-of-alberta-logo.png 1000w" sizes="(max-width: 268px) 100vw, 268px" /><br />
<a href="http://www.catolica.edu.sv/?page_id=3347"><img class="alignnone wp-image-3397" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-300x130.png" alt="uppsalalogo" width="258" height="112" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-300x130.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/uppsalalogo-1024x443.png 1024w" sizes="(max-width: 258px) 100vw, 258px" /></a><img class="alignnone wp-image-3398" src="http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen-300x150.png" alt="coop_externa-rrii_2016-02-26_becas_canada_elap_imagen" width="276" height="138" srcset="http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen-300x150.png 300w, http://www.catolica.edu.sv/wp-content/uploads/2016/01/coop_externa-rrii_2016-02-26_becas_canada_elap_imagen.png 600w" sizes="(max-width: 276px) 100vw, 276px" /></p>

		</div>
	</div>
</div></div></div></div></div><div class="container" ><div class="vc_row wpb_row vc_row-fluid mg-top-100 mg-bottom-100"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper">
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<div class="heading color-dark text-center mg-bottom-60">
<p><img class="alignnone size-full wp-image-4185" src="http://www.catolica.edu.sv/wp-content/uploads/2017/01/estrellas.jpg" alt="estrellas" width="56" height="25" /></p>
<h2 class="heading-color fs-38"><a style="color: #000000;" href="http://www.catolica.edu.sv/?post_type=tribe_events">Próximos eventos</a></h2>
</div>

		</div>
	</div>
                <div class="event style2  " >
                    <div data-plugin-options='{&quot;autoplay&quot;: true,&quot;loop&quot;:true,&quot;center&quot;:false,&quot;margin&quot;:0,&quot;animateOut&quot;:&quot;fadeOut&quot;,&quot;autoplayHoverPause&quot;:true,&quot;autoplayTimeout&quot;:5000,&quot;items&quot;:1,&quot;responsive&quot;:{},&quot;dots&quot;: true, &quot;nav&quot;:false}' class="owl-g5plus-shortcode owl-carousel">
                                                                            <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2018/01/slider-web-570x415.jpg" alt="Información para Graduación LX" title="Información para Graduación LX">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">enero 20 @ 8:00 am</span> - <span class="tribe-event-date-end">agosto 20 @ 5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=informacion-graduacion-lx" title="Información para Graduación LX" rel="bookmark">
                                                Información para Graduación LX                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">841</span>
                                                                                ENTREGA DE TOGAS, BIRRETE Y BORLAIndicaciones Serán entregadas ÚNICAMENTE del lunes 04 al sábado 09 de junio 2018, en horarios de 8:00 a.m. – 12:00 m. y de 3:00 – 7:00 p.m. en el primer nivel del edificio “C”. El sábado 09 de junio (Día del primer ensayo) ÚNICAMENTE se estará entregando de  9:00 a.m. [...]                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=informacion-graduacion-lx" title="Información para Graduación LX" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="" alt="Carreras semipresenciales bloque I" title="Carreras semipresenciales bloque I">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">febrero 3 @ 8:00 am</span> - <span class="tribe-event-date-end">abril 7 @ 8:20 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=carreras-semipresenciales-bloque-i" title="Carreras semipresenciales bloque I" rel="bookmark">
                                                Carreras semipresenciales bloque I                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">344</span>
                                                                                                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=carreras-semipresenciales-bloque-i" title="Carreras semipresenciales bloque I" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/SOLICITUD-DIFERIDOS-570x415.png" alt="Solicitud exámenes diferidos" title="Solicitud exámenes diferidos">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">marzo 19 @ 8:00 am</span> - <span class="tribe-event-date-end">marzo 24 @ 12:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=solicitud-examenes-diferidos" title="Solicitud exámenes diferidos" rel="bookmark">
                                                Solicitud exámenes diferidos                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">194</span>
                                                                                Según el artículo 20 del Reglamento de Evaluación del Rendimiento Académico Estudiantil, contemplado en el anuario académico: El estudiante que no se presente por causa justificada a una evaluación de fin de periodo podrá solicitar por escrito una evaluación diferida a Registro Académico. En el último período no habrá evaluación diferida. Y según el artículo [...]                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=solicitud-examenes-diferidos" title="Solicitud exámenes diferidos" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/DOC-GRADUACION-570x415.png" alt="Último día de entrega de documentos para graduación" title="Último día de entrega de documentos para graduación">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">marzo 20 @ 8:00 am</span> - <span class="tribe-event-time">6:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-entrega-de-documentos-para-graduacion" title="Último día de entrega de documentos para graduación" rel="bookmark">
                                                Último día de entrega de documentos para graduación                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">219</span>
                                                                                <p>Podrán ver todos los requisitos en: Registro Académico UNICAES Se solicita no dar credibilidad a la información que ofrezcan personas ajenas a Registro Académico en cuanto al registro de los títulos al MINED. Para obtener la solvencia económica deberá haber efectuado TODOS los pagos en Colecturía. Para mayor información pueden comunicarse al tel. 24840658 con  Rosalba [&hellip;]</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-entrega-de-documentos-para-graduacion" title="Último día de entrega de documentos para graduación" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="" alt="Cierre de instalaciones para actividades académicas" title="Cierre de instalaciones para actividades académicas">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">marzo 26 @ 8:00 am</span> - <span class="tribe-event-date-end">abril 2 @ 5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=cierre-de-instalaciones-para-actividades-academicas-2" title="Cierre de instalaciones para actividades académicas" rel="bookmark">
                                                Cierre de instalaciones para actividades académicas                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">2906</span>
                                                                                Recordatorio importante❗📢 ➡️ Se le recuerda a toda la comunidad universitaria que la UNICAES Sede Santa Ana y Facultad Multidisciplinaria de Ilobasco permanecerán cerradas por motivo de vacación colectiva, del 26 de marzo al 2 de abril. ➡️ No habrán actividades académicas ni administrativas, así como respuestas por diferentes medios (inbox, comentarios, llamadas y correos [...]                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=cierre-de-instalaciones-para-actividades-academicas-2" title="Cierre de instalaciones para actividades académicas" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/DIFERIDOS-570x415.png" alt="Exámenes diferidos" title="Exámenes diferidos">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">abril 3 @ 6:45 am</span> - <span class="tribe-event-date-end">abril 8 @ 8:20 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=examenes-diferidos-2" title="Exámenes diferidos" rel="bookmark">
                                                Exámenes diferidos                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">208</span>
                                                                                <p>Los horarios de realización están publicados en cada uno de los decanatos</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=examenes-diferidos-2" title="Exámenes diferidos" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/indexado-solo-pong-570x415.png" alt="Último día de pago de cuota" title="Último día de pago de cuota">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">abril 4 @ 8:00 am</span> - <span class="tribe-event-time">5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-pago-de-cuota-3" title="Último día de pago de cuota" rel="bookmark">
                                                Último día de pago de cuota                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">243</span>
                                                                                <p>Hoy es el último día para pagar cuota universitaria, en cualquier agencia del banco DAVIVIENDA y ventanilla en UNICAES, edificio &#8220;B&#8221; segundo nivel Horario de atención ventanilla UNICAES: 8:00 a.m. &#8211; 12:00 m. y de 1:00 &#8211; 5:00 p.m.</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-pago-de-cuota-3" title="Último día de pago de cuota" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/RETIRO-MATERIAS-570x415.png" alt="Último día para retirar materias" title="Último día para retirar materias">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">abril 9 @ 8:00 am</span> - <span class="tribe-event-time">5:30 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-para-retirar-materias" title="Último día para retirar materias" rel="bookmark">
                                                Último día para retirar materias                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">219</span>
                                                                                <p>Pasado este día ya no se podrá retirar materias. Puede encontrar el formulario aquí</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-para-retirar-materias" title="Último día para retirar materias" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/PARCIALES-570x415.png" alt="Exámenes parciales" title="Exámenes parciales">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">abril 30 @ 6:45 am</span> - <span class="tribe-event-date-end">mayo 5 @ 8:20 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=examenes-parciales-2" title="Exámenes parciales" rel="bookmark">
                                                Exámenes parciales                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">319</span>
                                                                                Hoy comienzan los exámenes parciales del segundo período del ciclo I-2018 Los horarios de parciales están publicados en cada uno de los decanatos ¡Bendiciones y muchos éxitos en sus parciales!                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=examenes-parciales-2" title="Exámenes parciales" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="" alt="Cierre de instalaciones para actividades académicas" title="Cierre de instalaciones para actividades académicas">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">mayo 1 @ 8:00 am</span> - <span class="tribe-event-time">6:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=cierre-de-instalaciones-para-actividades-academicas-9" title="Cierre de instalaciones para actividades académicas" rel="bookmark">
                                                Cierre de instalaciones para actividades académicas                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">230</span>
                                                                                "El trabajo más productivo es el que sale de las manos de un hombre contento" Victor Pauchet                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=cierre-de-instalaciones-para-actividades-academicas-9" title="Cierre de instalaciones para actividades académicas" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="" alt="Nuevo Ingreso Ciclo II-2018" title="Nuevo Ingreso Ciclo II-2018">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">mayo 2 @ 8:00 am</span> - <span class="tribe-event-date-end">junio 13 @ 5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=nuevo-ingreso-ciclo-ii-2018" title="Nuevo Ingreso Ciclo II-2018" rel="bookmark">
                                                Nuevo Ingreso Ciclo II-2018                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">192</span>
                                                                                Las inscripciones al Proceso de Ingreso para ciclo II 2018 están abiertas desde el 02 de mayo Inscríbete en línea También puedes venir a la UNICAES e inscribirte, solamente debes llenar la solicitud de inscripción del Proceso de Ingreso Ciclo II-2018 con tus datos personales y cancelar el costo total del Proceso de Ingreso de [...]                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=nuevo-ingreso-ciclo-ii-2018" title="Nuevo Ingreso Ciclo II-2018" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="" alt="Último día de pago de cuota" title="Último día de pago de cuota">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">mayo 4 @ 8:00 am</span> - <span class="tribe-event-time">5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-pago-de-cuota-5" title="Último día de pago de cuota" rel="bookmark">
                                                Último día de pago de cuota                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">99</span>
                                                                                <p>Hoy es el último día para pagar cuota universitaria, en cualquier agencia del banco DAVIVIENDA y ventanilla en UNICAES, edificio &#8220;B&#8221; segundo nivel Horario de atención ventanilla UNICAES: 8:00 a.m. &#8211; 12:00 m. y de 1:00 &#8211; 5:00 p.m.</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=ultimo-dia-de-pago-de-cuota-5" title="Último día de pago de cuota" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                    <div class="row-event-item">
                                <div class="col-md-6 col-sm-12 col-md-push-6 col-event-image">
                                    <img src="http://www.catolica.edu.sv/wp-content/uploads/2016/12/SOLICITUD-DIFERIDOS-570x415.png" alt="Solicitud de exámenes diferidos" title="Solicitud de exámenes diferidos">
                                </div>
                                <div class="col-md-6 col-sm-12 col-md-pull-6 col-event-content">
                                    <div class="content-middle-inner">
                                        <span class="tribe-event-date-start">mayo 7 @ 8:00 am</span> - <span class="tribe-event-date-end">mayo 12 @ 5:00 pm</span>                                        <h4>
                                            <a class="heading-color" href="http://www.catolica.edu.sv/?tribe_events=solicitud-de-examenes-diferidos-2" title="Solicitud de exámenes diferidos" rel="bookmark">
                                                Solicitud de exámenes diferidos                                            </a>
                                        </h4>
                                        <span class="event-comment">0</span>
                                                                                    <span class="event-view">228</span>
                                                                                <p>Según el artículo 20 del Reglamento de Evaluación del Rendimiento Académico Estudiantil, contemplado en el anuario académico: El estudiante que no se presente por causa justificada a una evaluación de fin de periodo podrá solicitar por escrito una evaluación diferida a Registro Académico. En el último período no habrá exaluación diferida. Y según el artículo [&hellip;]</p>
                                        <a class="bt bt-xs bt-bg bt-tertiary sm-mg-bottom-30" href="http://www.catolica.edu.sv/?tribe_events=solicitud-de-examenes-diferidos-2" title="Solicitud de exámenes diferidos" rel="bookmark">
                                            JOIN NOW                                        </a>
                                    </div>
                                </div>
                            </div>
                                                                    </div>
                </div>
            
	<div class="wpb_text_column wpb_content_element ">
		<div class="wpb_wrapper">
			<h5 style="text-align: center;"><a href="http://www.catolica.edu.sv/?post_type=tribe_events" target="_blank" rel="noopener noreferrer">(VER TODOS LOS EVENTOS)</a></h5>

		</div>
	</div>
</div></div></div></div></div><div class="fullwidth" ><div data-vc-parallax="1.5" data-overlay-color="rgba(136,12,10,1)" class="vc_row wpb_row vc_row-fluid vc_row-has-fill vc_row-o-equal-height vc_row-o-content-middle vc_row-flex vc_general vc_parallax vc_parallax-content-moving overlay-bg-vc-wapper"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper">                <div class="testimonial container style1 color-light pd-top-100 pd-bottom-100" >
                    <div class="fotorama" data-nav="thumbs" data-transition="crossfade" data-width="100%" data-height="240" data-autoplay="8000" data-thumbwidth="70" data-thumbheight="70" data-thumbmargin="10">
                                                    <div class="testimonial-item" data-thumb=" http://www.catolica.edu.sv/wp-content/uploads/2016/01/andrea-prueba.jpg">
                                <p>&quot;Estudiar en la UNICAES ha significado para mí conocer un nuevo mundo lleno de experiencias, donde se nos fortalece no solo el área profesional sino también el área de valores&quot;</p>
                                <h4 class="s-color">Andrea Ramos</h4>
                                <span>Estudiante de Licenciatura en Ciencias Jurídicas</span>
                            </div>
                                                        <div class="testimonial-item" data-thumb=" http://www.catolica.edu.sv/wp-content/uploads/2016/01/sayes-prueba.jpg">
                                <p>&quot;Como docente universitario una de mis mayores inspiraciones, ha sido el ver formados a los profesionales, y que luego se transforman en personas íntegras&quot;</p>
                                <h4 class="s-color">Lic. Carlos Sáyes</h4>
                                <span>Catedrático tiempo completo Facultad de Ciencias Empresariales</span>
                            </div>
                                                        <div class="testimonial-item" data-thumb=" http://www.catolica.edu.sv/wp-content/uploads/2016/01/Javier-Vanegas1.jpg">
                                <p>&quot;Consideré diversas universidades a nivel nacional y me fijé en la calidad, en la filosofía institucional y de cada profesional de UNICAES, por ese motivo decidí que quería estudiar aquí Ingeniería Industrial&quot;</p>
                                <h4 class="s-color">Ing. Javier Vanegas</h4>
                                <span>Ex alumno UNICAES</span>
                            </div>
                                                </div>
                </div>
            </div></div></div></div></div><div class="fullwidth" ><div class="vc_row wpb_row vc_row-fluid"><div class="wpb_column vc_column_container vc_col-sm-12"><div class="vc_column-inner "><div class="wpb_wrapper"><div class="vc_empty_space"  style="height: 100px" ><span class="vc_empty_space_inner"></span></div>
</div></div></div></div></div>
	</div>
	
</div>				</div>
                			</div>
								</main>			
			</div>
			<!-- Close Wrapper Content -->

			
							<footer  class="main-footer-wrapper dark">
					<div id="wrapper-footer">
						    <div class="footer-above-wrapper">
	    <div class="container">
		    <div class="footer-above-inner">
			    <div class="row">
				    					    <div class="col-md-6 sidebar">
						    <aside id="g5plus-footer-logo-3" class="widget widget-footer-logo">        <div class="footer-logo">
                            <a href="http://www.catolica.edu.sv"><img class="footer-logo-img" src="http://www.catolica.edu.sv/wp-content/uploads/2016/07/BLANCO-1.png" alt="UNICAES" /></a>
            	        	                </div>
        </aside>					    </div>
				    				    					    <div class="col-md-6 sidebar text-right">
						    <aside id="g5plus-social-profile-2" class="widget widget-social-profile"><ul class="social-profile s-rounded s-secondary s-md"><li><a title="Facebook" href="https://www.facebook.com/UNICAES/" target="_blank"><i class="fa fa-facebook"></i>Facebook</a></li>
<li><a title="Twitter" href="https://twitter.com/unicaes_sv/" target="_blank"><i class="fa fa-twitter"></i>Twitter</a></li>
<li><a title="Instagram" href="https://www.instagram.com/UNICAES_SV/" target="_blank"><i class="fa fa-instagram"></i>Instagram</a></li>
<li><a title="Youtube" href="https://www.youtube.com/channel/UCXDsbngj7qUa2wVlm9ogPvw" target="_blank"><i class="fa fa-youtube"></i>Youtube</a></li>
</ul></aside>					    </div>
				    			    </div>
		    </div>
	    </div>
    </div>
	<div class="main-footer">
		<div class="footer_inner clearfix">
	        <div class="footer_top_holder col-2">
	            <div class="container">
	                <div class="row footer-top-col-2 footer-7">
	                    <div class="sidebar footer-sidebar col-md-4 col-sm-12"><aside id="text-10" class="widget widget_text"><h4 class="widget-title">Nosotros</h4>			<div class="textwidget"><p style="text-align: justify;">La Universidad Católica de El Salvador tiene como Misión:
"La formación de personas, inspirada en los principios cristianos y en los conocimientos técnicos y científicos, orientada a una constante búsqueda de la verdad y del uso del saber, para contribuir a la tutela y desarrollo de la dignidad humana y de la sociedad, mediante la investigación, docencia y la proyección social."</p></div>
		</aside><aside id="text-11" class="widget widget_text"><h4 class="widget-title">contáctanos</h4>			<div class="textwidget"><ul class="footer-contact-us">
    <li>
        <i class="fa fa-map-marker"></i>
        <span>
            By pass carretera a Metapán y carretera Antigua hacia San Salvador.
        </span>
    </li>
   <li>
        <i class="fa fa-phone"></i>
        <span>
            2484-0600
            Fax 2441-2655
        </span>
    </li>
    <li>
        <i class="fa fa-envelope"></i>
        <span>
            catolica@catolica.edu.sv
        </span>
    </li>
    
</ul></div>
		</aside></div><div class="sidebar footer-sidebar col-md-8 col-sm-12"><aside id="search-4" class="widget widget_search"><h4 class="widget-title">Búsqueda</h4><form class="search-form" method="get" id="searchform" action="http://www.catolica.edu.sv/">
                <input type="text" value="" name="s" id="s"  placeholder="INTRODUZCA PALABRA">
                <button type="submit"><i class="fa fa-search"></i>Search</button>
     		</form></aside><aside id="null-instagram-feed-3" class="widget null-instagram-feed"><h4 class="widget-title">Instagram</h4>Instagram has returned invalid data.<p class="clear"><a href="//instagram.com/unicaes_sv/" rel="me" target="_self" class="">Síguenos</a></p></aside><aside id="text-17" class="widget widget_text"><h4 class="widget-title">Visitantes</h4>			<div class="textwidget"><script type="text/javascript" id="clustrmaps" src="//cdn.clustrmaps.com/map_v2.js?d=lyWFEbmgCk5R_I5Zj1qswU_Y6c_OKFRCisH0apVT8Q0&cl=ffffff&w=a"></script></div>
		</aside></div>	                </div>
	            </div>
	        </div>
		</div>
	</div>
	<div class="bottom-bar-wrapper">
		<div class="container">
			<div class="bottom-bar-inner">
				<div class="row">
											<div class="col-md-6 sidebar text-left">
							<aside id="nav_menu-2" class="dark widget widget_nav_menu"><div class="menu-footer-menu-container"><ul id="menu-footer-menu" class="menu"><li id="menu-item-889" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-home current-menu-item page_item page-item-321 current_page_item menu-item-889"><a href="http://www.catolica.edu.sv/">INICIO</a></li>
<li id="menu-item-2073" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-2073"><a href="http://www.catolica.edu.sv/?page_id=1057">Oferta Académica</a></li>
<li id="menu-item-2074" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-2074"><a href="http://www.catolica.edu.sv/?page_id=671">Postgrado</a></li>
<li id="menu-item-899" class="menu-item menu-item-type-post_type menu-item-object-page menu-item-899"><a href="http://www.catolica.edu.sv/?page_id=861">Noticias</a></li>
</ul></div></aside>						</div>
																<div class="col-md-6 sidebar text-right">
							<aside id="text-4" class="dark widget widget_text">			<div class="textwidget">UNIVERSIDAD CATÓLICA DE EL SALVADOR</div>
		</aside>						</div>
									</div>
			</div>
		</div>
	</div>
					</div>
				</footer>
					</div>
		<!-- Close Wrapper -->

			<!-- analytics-code google analytics tracking code --><script>
	(function(i,s,o,g,r,a,m){i['GoogleAnalyticsObject']=r;i[r]=i[r]||function(){
			(i[r].q=i[r].q||[]).push(arguments)},i[r].l=1*new Date();a=s.createElement(o),
		m=s.getElementsByTagName(o)[0];a.async=1;a.src=g;m.parentNode.insertBefore(a,m)
	})(window,document,'script','//www.google-analytics.com/analytics.js','ga');

	ga('create', 'UA-96475387-1', 'auto');
	ga('send', 'pageview');

</script><!--  -->		<script>
		( function ( body ) {
			'use strict';
			body.className = body.className.replace( /\btribe-no-js\b/, 'tribe-js' );
		} )( document.body );
		</script>
		<script type="text/javascript">                                    </script><script type='text/javascript'> /* <![CDATA[ */var tribe_l10n_datatables = {"aria":{"sort_ascending":": activate to sort column ascending","sort_descending":": activate to sort column descending"},"length_menu":"Show _MENU_ entries","empty_table":"No data available in table","info":"Showing _START_ to _END_ of _TOTAL_ entries","info_empty":"Showing 0 to 0 of 0 entries","info_filtered":"(filtered from _MAX_ total entries)","zero_records":"No matching records found","search":"Search:","all_selected_text":"All items on this page were selected. ","select_all_link":"Select all pages","clear_selection":"Clear Selection.","pagination":{"all":"All","next":"Siguiente","previous":"Previous"},"select":{"rows":{"0":"","_":": Selected %d rows","1":": Selected 1 row"}},"datepicker":{"dayNames":["domingo","lunes","martes","mi\u00e9rcoles","jueves","viernes","s\u00e1bado"],"dayNamesShort":["Dom","Lun","Mar","Mie","Jue","Vie","Sab"],"dayNamesMin":["D","L","M","X","J","V","S"],"monthNames":["enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre"],"monthNamesShort":["enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre"],"nextText":"Siguiente","prevText":"Anterior","currentText":"Hoy","closeText":"Hecho"}};/* ]]> */ </script><link rel='stylesheet' property='stylesheet' id='rs-icon-set-fa-icon-css'  href='http://www.catolica.edu.sv/wp-content/plugins/revslider/public/assets/fonts/font-awesome/css/font-awesome.css' type='text/css' media='all' />		<script type="text/javascript">
			function revslider_showDoubleJqueryError(sliderID) {
				var errorMessage = "Revolution Slider Error: You have some jquery.js library include that comes after the revolution files js include.";
				errorMessage += "<br> This includes make eliminates the revolution slider libraries, and make it not work.";
				errorMessage += "<br><br> To fix it you can:<br>&nbsp;&nbsp;&nbsp; 1. In the Slider Settings -> Troubleshooting set option:  <strong><b>Put JS Includes To Body</b></strong> option to true.";
				errorMessage += "<br>&nbsp;&nbsp;&nbsp; 2. Find the double jquery.js include and remove it.";
				errorMessage = "<span style='font-size:16px;color:#BC0C06;'>" + errorMessage + "</span>";
					jQuery(sliderID).show().html(errorMessage);
			}
		</script>
				<script type="text/javascript">
			function revslider_showDoubleJqueryError(sliderID) {
				var errorMessage = "Revolution Slider Error: You have some jquery.js library include that comes after the revolution files js include.";
				errorMessage += "<br> This includes make eliminates the revolution slider libraries, and make it not work.";
				errorMessage += "<br><br> To fix it you can:<br>&nbsp;&nbsp;&nbsp; 1. In the Slider Settings -> Troubleshooting set option:  <strong><b>Put JS Includes To Body</b></strong> option to true.";
				errorMessage += "<br>&nbsp;&nbsp;&nbsp; 2. Find the double jquery.js include and remove it.";
				errorMessage = "<span style='font-size:16px;color:#BC0C06;'>" + errorMessage + "</span>";
					jQuery(sliderID).show().html(errorMessage);
			}
		</script>
		<link rel='stylesheet' id='g5plus_vc_extend_css-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/themes/academia/assets/vc-extend/css/vc-customize.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='flexslider-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/flexslider/flexslider.min.css?ver=4.11.2.1' type='text/css' media='all' />
<link rel='stylesheet' id='academia_event_css-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/academia-framework/includes/shortcodes/event/assets/css/event.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='vc_google_fonts_abril_fatfaceregular-css'  property='stylesheet' href='//fonts.googleapis.com/css?family=Abril+Fatface%3Aregular&#038;subset=latin&#038;ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='academia_testimonial_css-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/academia-framework/includes/shortcodes/testimonial/assets/css/testimonial.min.css?ver=4.7.9' type='text/css' media='all' />
<link rel='stylesheet' id='academia_fotorama_css-css'  property='stylesheet' href='http://www.catolica.edu.sv/wp-content/plugins/academia-framework/includes/shortcodes/testimonial/assets/css/fotorama.css?ver=4.7.9' type='text/css' media='all' />
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/contact-form-7/includes/js/jquery.form.min.js?ver=3.51.0-2014.06.20'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var _wpcf7 = {"recaptcha":{"messages":{"empty":"Por favor, prueba que no eres un robot."}},"cached":"1"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/contact-form-7/includes/js/scripts.js?ver=4.7'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/bootstrap/js/bootstrap.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/js/plugin.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/smoothscroll/SmoothScroll.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/jquery.jPlayer/jquery.jplayer.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/plugins/slick/js/slick.min.js?ver=4.7.9'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var g5plus_framework_ajax_url = "http:\/\/www.catolica.edu.sv\/wp-admin\/admin-ajax.php?activate-multi=true";
var g5plus_framework_theme_url = "http:\/\/www.catolica.edu.sv\/wp-content\/themes\/academia\/";
var g5plus_framework_site_url = "http:\/\/www.catolica.edu.sv";
/* ]]> */
</script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/js/main.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-includes/js/wp-embed.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/js/dist/js_composer_front.min.js?ver=4.11.2.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/assets/vc-extend/js/vc_extend.min.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/flexslider/jquery.flexslider-min.js?ver=4.11.2.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/vc_accordion/vc-accordion.min.js?ver=4.11.2.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/vc-tta-autoplay/vc-tta-autoplay.min.js?ver=4.11.2.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/js_composer/assets/lib/bower/skrollr/dist/skrollr.min.js?ver=4.11.2.1'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/plugins/academia-framework/includes/shortcodes/testimonial/assets/js/fotorama.js?ver=4.7.9'></script>
<script type='text/javascript' src='http://www.catolica.edu.sv/wp-content/themes/academia/g5plus-framework/xmenu/assets/js/app.min.js?ver=1.0.0.0'></script>
<script>jQuery("style#g5plus_custom_style").append("@media screen and (min-width: 992px) {}");</script><script>jQuery("style#g5plus_custom_style").append("@media screen and (min-width: 992px) {}");</script></body>
</html> <!-- end of site. what a ride! -->
<!-- Performance optimized by W3 Total Cache. Learn more: https://www.w3-edge.com/products/

 Served from: www.catolica.edu.sv @ 2018-03-19 22:02:38 by W3 Total Cache -->