<!DOCTYPE html>
<!--[if lt IE 7]>      <html class="no-js lt-ie9 lt-ie8 lt-ie7" lang="es-ES"> <![endif]-->
<!--[if IE 7]>         <html class="no-js lt-ie9 lt-ie8" lang="es-ES"> <![endif]-->
<!--[if IE 8]>         <html class="no-js lt-ie9" lang="es-ES"> <![endif]-->
<!--[if gt IE 8]><!--> <html class="no-js" lang="es-ES"> <!--<![endif]-->
	<head>
		<title>MINSAL | Sitio Oficial del Ministerio de Salud de El Salvador</title>
		
		<!-- Default Meta Tags -->
		<meta charset="UTF-8">

<link href="//www.google-analytics.com" rel="dns-prefetch">

<meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">

<meta name="viewport" content="width=device-width,initial-scale=1.0,user-scalable=yes">

<meta name="keywords" content="El Salvador, Ministerio, Salud, Convocatorias de Prensa, Servicios, Estadísticas, Adjudicaciones y Contrataciones, Programas de Salud, Vigilancia Epidemiológica, Guía de Servicios, Actividades de Titulares" />

<meta name="description" content="Sitio Oficial del Ministerio de Salud de El Salvador">
<link rel="shortcut icon" href="http://www.salud.gob.sv/wp-content/uploads/2015/01/favicon.png">		




<link rel="pingback" href="http://www.salud.gob.sv/xmlrpc.php" />

		<!-- Facebook integration -->
  

<meta property="og:site_name" content="MINSAL">

<meta property="og:url" content="http://www.salud.gob.sv"/>  
<meta property="og:type" content="website" />
<meta property="og:title" content="MINSAL  Sitio Oficial del Ministerio de Salud de El Salvador">
<meta property="og:description" content="Sitio Oficial del Ministerio de Salud de El Salvador">



		<!-- css + javascript -->
		<link rel='dns-prefetch' href='//ajax.googleapis.com' />
<link rel='dns-prefetch' href='//s.w.org' />
<link rel="alternate" type="application/rss+xml" title="MINSAL &raquo; Feed" href="http://www.salud.gob.sv/feed/" />
<link rel="alternate" type="application/rss+xml" title="MINSAL &raquo; RSS de los comentarios" href="http://www.salud.gob.sv/comments/feed/" />
<link rel="alternate" type="text/calendar" title="MINSAL &raquo; iCal Feed" href="http://www.salud.gob.sv/events/?ical=1" />
<link rel="alternate" type="application/rss+xml" title="MINSAL &raquo; Inicio RSS de los comentarios" href="http://www.salud.gob.sv/inicio-2/feed/" />
		<script type="text/javascript">
			window._wpemojiSettings = {"baseUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/72x72\/","ext":".png","svgUrl":"https:\/\/s.w.org\/images\/core\/emoji\/2.4\/svg\/","svgExt":".svg","source":{"concatemoji":"http:\/\/www.salud.gob.sv\/wp-includes\/js\/wp-emoji-release.min.js?ver=4.9.4"}};
			!function(a,b,c){function d(a,b){var c=String.fromCharCode;l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,a),0,0);var d=k.toDataURL();l.clearRect(0,0,k.width,k.height),l.fillText(c.apply(this,b),0,0);var e=k.toDataURL();return d===e}function e(a){var b;if(!l||!l.fillText)return!1;switch(l.textBaseline="top",l.font="600 32px Arial",a){case"flag":return!(b=d([55356,56826,55356,56819],[55356,56826,8203,55356,56819]))&&(b=d([55356,57332,56128,56423,56128,56418,56128,56421,56128,56430,56128,56423,56128,56447],[55356,57332,8203,56128,56423,8203,56128,56418,8203,56128,56421,8203,56128,56430,8203,56128,56423,8203,56128,56447]),!b);case"emoji":return b=d([55357,56692,8205,9792,65039],[55357,56692,8203,9792,65039]),!b}return!1}function f(a){var c=b.createElement("script");c.src=a,c.defer=c.type="text/javascript",b.getElementsByTagName("head")[0].appendChild(c)}var g,h,i,j,k=b.createElement("canvas"),l=k.getContext&&k.getContext("2d");for(j=Array("flag","emoji"),c.supports={everything:!0,everythingExceptFlag:!0},i=0;i<j.length;i++)c.supports[j[i]]=e(j[i]),c.supports.everything=c.supports.everything&&c.supports[j[i]],"flag"!==j[i]&&(c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&c.supports[j[i]]);c.supports.everythingExceptFlag=c.supports.everythingExceptFlag&&!c.supports.flag,c.DOMReady=!1,c.readyCallback=function(){c.DOMReady=!0},c.supports.everything||(h=function(){c.readyCallback()},b.addEventListener?(b.addEventListener("DOMContentLoaded",h,!1),a.addEventListener("load",h,!1)):(a.attachEvent("onload",h),b.attachEvent("onreadystatechange",function(){"complete"===b.readyState&&c.readyCallback()})),g=c.source||{},g.concatemoji?f(g.concatemoji):g.wpemoji&&g.twemoji&&(f(g.twemoji),f(g.wpemoji)))}(window,document,window._wpemojiSettings);
		</script>
		<style type="text/css">
img.wp-smiley,
img.emoji {
	display: inline !important;
	border: none !important;
	box-shadow: none !important;
	height: 1em !important;
	width: 1em !important;
	margin: 0 .07em !important;
	vertical-align: -0.1em !important;
	background: none !important;
	padding: 0 !important;
}
</style>
<link rel='stylesheet' id='google-language-translator-css'  href='http://www.salud.gob.sv/wp-content/plugins/google-language-translator/css/style.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='bootstrap_tab-css'  href='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/css/bootstrap_tab.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='bootstrap_dropdown-css'  href='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/css/bootstrap_dropdown.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='ert_tab_icon_css-css'  href='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/css/res_tab_icon.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='contact-form-7-css'  href='http://www.salud.gob.sv/wp-content/plugins/contact-form-7/includes/css/styles.css?ver=5.0' type='text/css' media='all' />
<link rel='stylesheet' id='jquery-ui-theme-css'  href='http://ajax.googleapis.com/ajax/libs/jqueryui/1.11.4/themes/humanity/jquery-ui.min.css?ver=1.11.4' type='text/css' media='all' />
<link rel='stylesheet' id='jquery-ui-timepicker-css'  href='http://www.salud.gob.sv/wp-content/plugins/contact-form-7-datepicker/js/jquery-ui-timepicker/jquery-ui-timepicker-addon.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='font-awesome-css'  href='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/font-awesome/css/font-awesome.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='wpdm-bootstrap-css'  href='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/bootstrap/css/bootstrap.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='wpdm-front-css'  href='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/css/front.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='showbiz-settings-css'  href='http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/css/settings.css?ver=1.7.2' type='text/css' media='all' />
<link rel='stylesheet' id='fancybox-css'  href='http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/fancybox/jquery.fancybox.css?ver=1.7.2' type='text/css' media='all' />
<link rel='stylesheet' id='wk-styles-css'  href='http://www.salud.gob.sv/wp-content/plugins/widgetkit/cache/wk-styles-d5b6099f.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='wordpress-popular-posts-css-css'  href='http://www.salud.gob.sv/wp-content/plugins/wordpress-popular-posts/public/css/wpp.css?ver=4.0.13' type='text/css' media='all' />
<link rel='stylesheet' id='chosen-css'  href='http://www.salud.gob.sv/wp-content/plugins/wp-job-manager/assets/css/chosen.css?ver=1.1.0' type='text/css' media='all' />
<link rel='stylesheet' id='wp-job-manager-frontend-css'  href='http://www.salud.gob.sv/wp-content/plugins/wp-job-manager/assets/css/frontend.css?ver=1.29.3' type='text/css' media='all' />
<link rel='stylesheet' id='rokbox.css-css'  href='http://www.salud.gob.sv/wp-content/plugins/wp_rokbox/assets/styles/rokbox.css?ver=2.50.5' type='text/css' media='all' />
<link rel='stylesheet' id='dashicons-css'  href='http://www.salud.gob.sv/wp-includes/css/dashicons.min.css?ver=4.9.4' type='text/css' media='all' />
<link rel='stylesheet' id='spu-public-css-css'  href='http://www.salud.gob.sv/wp-content/plugins/popups/public/assets/css/public.css?ver=1.9.1.1' type='text/css' media='all' />
<link rel='stylesheet' id='tablepress-default-css'  href='http://www.salud.gob.sv/wp-content/plugins/tablepress/css/default.min.css?ver=1.9' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-flexslider-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/flexslider/flexslider-custom.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-icon-social-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/font-icons/social-icons/css/zocial.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-icon-entypo-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/font-icons/entypo/css/entypo.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-icon-symbol-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/font-icons/symbol/css/symbol.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-swipebox-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/swipebox/swipebox.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-bootstrap-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/bootstrap/css/bootstrap.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='vwcss-theme-css'  href='http://www.salud.gob.sv/wp-content/themes/RedSV/css/theme.css?ver=1.9.0' type='text/css' media='all' />
<link rel='stylesheet' id='pcs-styles-css'  href='http://www.salud.gob.sv/wp-content/plugins/post-content-shortcodes/styles/default-styles.css?ver=1.0' type='text/css' media='screen' />
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/jquery.js?ver=1.12.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/jquery-migrate.min.js?ver=1.4.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/google-language-translator/js/load-flags.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/wp_rokbox/assets/js/mootools.js?ver=1.4.5'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/bootstrap/js/bootstrap.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/js/front.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/js/chosen.jquery.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/fancybox/jquery.fancybox.pack.js?ver=1.7.2'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/js/jquery.themepunch.tools.min.js?ver=1.7.2'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/js/jquery.themepunch.showbizpro.min.js?ver=1.7.2'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/widgetkit/cache/uikit-3e16fcfd.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/widgetkit/cache/wk-scripts-9dccfd4a.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/wp-featured-content-slider/scripts/jquery.cycle.all.2.72.js?ver=1.3'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/wp_rokbox/assets/js/rokbox.js?ver=2.50.5'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var instant_search = {"blog_url":"http:\/\/www.salud.gob.sv","ajax_url":"http:\/\/www.salud.gob.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/instant-search/instant-search.js?ver=4.9.4'></script>
<meta name="generator" content="WordPress Download Manager 2.9.69" />
<link rel='https://api.w.org/' href='http://www.salud.gob.sv/wp-json/' />
<link rel="EditURI" type="application/rsd+xml" title="RSD" href="http://www.salud.gob.sv/xmlrpc.php?rsd" />
<link rel="wlwmanifest" type="application/wlwmanifest+xml" href="http://www.salud.gob.sv/wp-includes/wlwmanifest.xml" /> 
<link rel="canonical" href="http://www.salud.gob.sv/" />
<link rel='shortlink' href='http://www.salud.gob.sv/' />
<link rel="alternate" type="application/json+oembed" href="http://www.salud.gob.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fwww.salud.gob.sv%2F" />
<link rel="alternate" type="text/xml+oembed" href="http://www.salud.gob.sv/wp-json/oembed/1.0/embed?url=http%3A%2F%2Fwww.salud.gob.sv%2F&#038;format=xml" />
<meta name="framework" content="Alkivia Framework 0.8" />
<script type='text/javascript'>
/* <![CDATA[ */
// Comprehensive Google Map plugin v9.1.2
var CGMPGlobal = {"ajaxurl":"http:\/\/www.salud.gob.sv\/wp-admin\/admin-ajax.php","noBubbleDescriptionProvided":"No description provided","geoValidationClientRevalidate":"REVALIDATE","cssHref":"http:\/\/www.salud.gob.sv\/wp-content\/plugins\/comprehensive-google-map-plugin\/style.css?ver=9.1.2","language":"en","customMarkersUri":"http:\/\/www.salud.gob.sv\/wp-content\/plugins\/comprehensive-google-map-plugin\/assets\/css\/images\/markers\/","kml":"[TITLE] [MSG] ([STATUS])","kmlDocInvalid":"The KML file is not a valid KML, KMZ or GeoRSS document.","kmlFetchError":"The KML file could not be fetched.","kmlLimits":"The KML file exceeds the feature limits of KmlLayer.","kmlNotFound":"The KML file could not be found. Most likely it is an invalid URL, or the document is not publicly available.","kmlRequestInvalid":"The KmlLayer is invalid.","kmlTimedOut":"The KML file could not be loaded within a reasonable amount of time.","kmlTooLarge":"The KML file exceeds the file size limits of KmlLayer.","kmlUnknown":"The KML file failed to load for an unknown reason.","address":"Address","streetView":"Street View","directions":"Directions","toHere":"To here","fromHere":"From here","mapFillViewport":"true","timestamp":"094536421d","ajaxCacheMapAction":"cgmp_ajax_cache_map_action","sep":"{}"}
/* ]]> */
</script>

        <script>
            var wpdm_site_url = 'http://www.salud.gob.sv/';
            var wpdm_home_url = 'http://www.salud.gob.sv/';
            var ajax_url = 'http://www.salud.gob.sv/wp-admin/admin-ajax.php';
            var wpdm_ajax_url = 'http://www.salud.gob.sv/wp-admin/admin-ajax.php';
            var wpdm_ajax_popup = '0';
        </script>


        <style type="text/css">#google_language_translator a {display: none !important; }.goog-te-gadget {color:transparent !important;}.goog-te-gadget { font-size:0px !important; }.goog-branding { display:none; }.goog-tooltip {display: none !important;}.goog-tooltip:hover {display: none !important;}.goog-text-highlight {background-color: transparent !important; border: none !important; box-shadow: none !important;}#flags { display:none; }#google_language_translator {color: transparent;}body { top:0px !important; }</style><link rel="stylesheet" href="http://www.salud.gob.sv/wp-content/plugins/multi-column-taxonomy-list/css/multi-column-taxonomy-link.css" type="text/css" />    <style type="text/css" media="screen">
      div.printfriendly a, div.printfriendly a:link, div.printfriendly a:hover, div.printfriendly a:visited {
        text-decoration: none;
        border: none;
      }
    </style>
   
<style>
.scroll-back-to-top-wrapper {
    position: fixed;
	opacity: 0;
	visibility: hidden;
	overflow: hidden;
	text-align: center;
	z-index: 99999999;
    background-color: #1e73be;
	color: #eeeeee;
	width: 50px;
	height: 48px;
	line-height: 48px;
	right: 30px;
	bottom: 30px;
	padding-top: 2px;
	border-top-left-radius: 10px;
	border-top-right-radius: 10px;
	border-bottom-right-radius: 10px;
	border-bottom-left-radius: 10px;
	-webkit-transition: all 0.5s ease-in-out;
	-moz-transition: all 0.5s ease-in-out;
	-ms-transition: all 0.5s ease-in-out;
	-o-transition: all 0.5s ease-in-out;
	transition: all 0.5s ease-in-out;
}
.scroll-back-to-top-wrapper:hover {
	background-color: #7499bf;
  color: #eeeeee;
}
.scroll-back-to-top-wrapper.show {
    visibility:visible;
    cursor:pointer;
	opacity: 1.0;
}
.scroll-back-to-top-wrapper i.fa {
	line-height: inherit;
}
.scroll-back-to-top-wrapper .fa-lg {
	vertical-align: 0;
}
</style><script type="text/javascript">if (typeof RokBoxSettings == 'undefined') RokBoxSettings = {pc: '100'};</script>
<script type="text/javascript" src="http://www.salud.gob.sv/wp-content/plugins/zd-youtube-flv-player/js/swfobject.js"></script>
<meta name="tec-api-version" content="v1"><meta name="tec-api-origin" content="http://www.salud.gob.sv"><link rel="https://theeventscalendar.com/" href="http://www.salud.gob.sv/wp-json/tribe/events/v1/" />	<style type="text/css" id="custom-background-css">
	body.custom-background.site-layout-boxed
	, body.custom-background.site-layout-full-large #off-canvas-body-inner
	, body.custom-background.site-layout-full-medium #off-canvas-body-inner
	{ background-color: #d6eaf8; }
	</style>
	<link href='http://fonts.googleapis.com/css?family=Roboto:400,400italic,700,700italic,700,700italic|Open+Sans:400,400italic,700,700italic,400,400italic&#038;subset=latin,latin-ext,cyrillic,cyrillic-ext,greek-ext,greek,vietnamese' rel='stylesheet' type='text/css'>	<style type="text/css">
				
				
		::selection { color: white; background-color: #3facd6; }
		h1, h2, h3, h4, h5, h6 {
			font-family: Roboto, sans-serif;
			font-weight: 700;
			color: #000000;
		}
		h1 { line-height: 1.1; }
		h2 { line-height: 1.2; }
		h3, h4, h5, h6 { line-height: 1.4; }
		body {
			font-family: Open Sans, sans-serif;
			font-size: 14px;
			font-weight: 400;
			color: #545454;
		}

		.header-font,
		woocommerce div.product .woocommerce-tabs ul.tabs li, .woocommerce-page div.product .woocommerce-tabs ul.tabs li, .woocommerce #content div.product .woocommerce-tabs ul.tabs li, .woocommerce-page #content div.product .woocommerce-tabs ul.tabs li
		{ font-family: Roboto, sans-serif; font-weight: 700; }
		.header-font-color { color: #000000; }

		.wp-caption p.wp-caption-text {
			color: #000000;
			border-bottom-color: #000000;
		}
		
		.body-font { font-family: Open Sans, sans-serif; font-weight: 400; }

		/* Only header font, No font-weight */
		.mobile-nav,
		.top-nav,
		.comment .author > span, .pingback .author > span, 
		.label, .tagcloud a,
		.woocommerce .product_meta .post-tags a,
		.bbp-topic-tags a,
		.woocommerce div.product span.price, .woocommerce-page div.product span.price, .woocommerce #content div.product span.price, .woocommerce-page #content div.product span.price, .woocommerce div.product p.price, .woocommerce-page div.product p.price, .woocommerce #content div.product p.price, .woocommerce-page #content div.product p.price,
		.main-nav .menu-link { font-family: Roboto, sans-serif; }

		/* Primary Color */
		.primary-bg,
		.label, .tagcloud a,
		.woocommerce nav.woocommerce-pagination ul li span.current, .woocommerce-page nav.woocommerce-pagination ul li span.current, .woocommerce #content nav.woocommerce-pagination ul li span.current, .woocommerce-page #content nav.woocommerce-pagination ul li span.current, .woocommerce nav.woocommerce-pagination ul li a:hover, .woocommerce-page nav.woocommerce-pagination ul li a:hover, .woocommerce #content nav.woocommerce-pagination ul li a:hover, .woocommerce-page #content nav.woocommerce-pagination ul li a:hover, .woocommerce nav.woocommerce-pagination ul li a:focus, .woocommerce-page nav.woocommerce-pagination ul li a:focus, .woocommerce #content nav.woocommerce-pagination ul li a:focus, .woocommerce-page #content nav.woocommerce-pagination ul li a:focus,
		#pagination > span {
			background-color: #3facd6;
		}
		a, .social-share a:hover, .site-social-icons a:hover,
		.bbp-topic-header a:hover,
		.bbp-forum-header a:hover,
		.bbp-reply-header a:hover { color: #3facd6; }
		.button-primary { color: #3facd6; border-color: #3facd6; }
		.primary-border { border-color: #3facd6; }

		/* Top-bar Colors */
		.top-bar {
			background-color: #023f62;
			color: #ffffff;
		}

		#open-mobile-nav, .top-nav  a, .top-bar-right > a {
			color: #ffffff;
		}

		#open-mobile-nav:hover, .top-nav  a:hover, .top-bar-right > a:hover {
			background-color: #3facd6;
			color: #ffffff;
		}

		.top-nav .menu-item:hover { background-color: #3facd6; }
		.top-nav .menu-item:hover > a { color: #ffffff; }

		/* Header Colors */
		.main-bar {
			background-color: #0368a1;
			color: #ffffff;
		}

		/* Main Navigation Colors */
		.main-nav-bar {
			background-color: #023f62;
		}

		.main-nav-bar, .main-nav > .menu-item > a {
			color: #ffffff;
		}

		.main-nav .menu-item:hover > .menu-link,
		.main-nav > .current-menu-ancestor > a,
		.main-nav > .current-menu-item > a {
			background-color: #3facd6;
			color: #ffffff;
		}

		/* Widgets */
		.widget_vw_widget_social_subscription .social-subscription:hover .social-subscription-icon { background-color: #3facd6; }
		.widget_vw_widget_social_subscription .social-subscription:hover .social-subscription-count { color: #3facd6; }

		.widget_vw_widget_categories a:hover { color: #3facd6; }

		/* Footer Colors */
		#footer {
			background-color: #045583;
		}

		#footer .widget-title {
			color: #3facd6;
		}

		#footer,
		#footer .title,
		#footer .comment-author,
		#footer .social-subscription-count
		{ color: #ffffff; }

		.copyright {
			background-color: #045583;
		}
		.copyright, .copyright a {
			color: #ffffff;
		}

		/* Custom Styles */
				/* TABLA CONGRESO INT REFORMA DE LA SALUD 2017*/
table.congreso {font-size:12px;color:#333333;width:100%;border-width: 1px;border-color: #729ea5;border-collapse: collapse;}
table.congreso th {font-size:12px;background-color:#00AFEF;border-width: 1px;padding: 8px;border-style: solid;border-color: #729ea5;text-align:center;}
/*table.congreso tr {background-color:#d4e3e5;}*/
table.congreso td {font-size:12px;border-width: 1px;padding: 8px;border-style: solid;border-color: #729ea5;}


.img2016 {
display: block;
margin: auto;
width: 40%;
}

/* Menu UISP-2016 */
.menu_post 1{
    background-color: #006699;
    border: none;
    color: white;
    padding: 8px 8px;
    text-align: center;
    text-decoration: none;
    display: inline-block;
    font-size: 10px;
    cursor: pointer;
    float: center;
}

.menu_post1:hover {
    background-color: #FFFFFF;
}

.button {
    background-color: #f4511e; /* Green */
    border: none;
    border-radius: 4px;
    color: white;
    padding: 15px 25px;
    text-align: center;
    text-decoration: none;
    display: inline-block;
    font-size: 10px;
    cursor: pointer;
    float: right;
}

.button:hover {
    background-color:  #b3b6b7 ;
}

.menu_post {
    background-color: #006699; /* Green */
    border: none;
    color: white;
    padding: 10px 8px;
    text-align: center;
    text-decoration: none;
    display: inline-block;
    font-size: 10px;
    cursor: pointer;
    float: center;
}

.menu_post:hover {
    background-color: #6699CC;
}



.main-nav > .menu-item > .menu-link {
    font-size: 16px;
}

/*MENU Y SUBMENUS EN NEGRILLA*/
.main-nav-bar, .main-nav > .menu-item > a {
    font-weight:bold !important;
}


/* Mostrar subniveles del menu */
/*Cambiar valor header.php line 128 depth' => 0, estaba:2 y quedo 0*/
nav ul ul ul {
   
  position: absolute;
    margin-top: -38px;
    left:100%;
      min-width:325px;
}

table.tftable {font-size:12px;color:#333333;width:100%;border-width: 1px;border-color: #729ea5;border-collapse: collapse;}
table.tftable th {font-size:12px;background-color:#acc8cc;border-width: 1px;padding: 8px;border-style: solid;border-color: #729ea5;text-align:center;}
table.tftable tr {background-color:#d4e3e5;}
table.tftable td {font-size:12px;border-width: 1px;padding: 8px;border-style: solid;border-color: #729ea5;}

/* Estilo del div para el boton de logout */
#estilo1{color:#FFFFFF;background:orange;}

.su-spoiler.my-custom-spoiler {}
.su-spoiler.my-custom-spoiler .su-spoiler-title { background-color: #6699CC }
.su-spoiler.my-custom-spoiler .su-spoiler-title .su-spoiler-icon,
.su-spoiler.su-spoiler-closed.my-custom-spoiler .su-spoiler-title .su-spoiler-icon {
left: 3px;
background-color: #fff;
}
.su-spoiler.my-custom-spoiler .su-spoiler-content { background-color: #eeeeee }
.su-spoiler-title {color: #000000}
#box
{
    height: 34px;
    width: 700px;
    background: #073763;
    font-size: 20px;
    font-style: "Roboto", sans-serif;
    color: #FFF;
    text-align: center;
    margin-top: 0px;
    margin-left: 5px;
    font-weight: bold;
    vertical-align: middle;
    display: table-cell;
    border-radius: 5px;
}


.su-spoiler.my-custom-spoiler {}
.su-spoiler.my-custom-spoiler .su-spoiler-title { background-color: #6699CC }
.su-spoiler.my-custom-spoiler .su-spoiler-title .su-spoiler-icon,
.su-spoiler.su-spoiler-closed.my-custom-spoiler .su-spoiler-title .su-spoiler-icon {
left: 3px;
background-color: #fff;
}
.su-spoiler.my-custom-spoiler .su-spoiler-content { background-color: #eeeeee }
.su-spoiler-title {color: #000000}
#box1
{
    height: 50px;
    line-height: 50px;
    width: 380px;
    background: #073763;
    font-size: 130%;
    font-style: "Roboto", sans-serif;
    color: #FFF;
    text-align: center;
    margin-top: 0px;
    margin-left: 5px;
    font-weight: bold;
    vertical-align: middle;
    display: block;
    float: left;
    border-radius: 5px;
    padding: 0px 0px 0px 0px;
    margin-bottom: 5px; 
    position: relative;
}


.su-spoiler.my-custom-spoiler {}
.su-spoiler.my-custom-spoiler .su-spoiler-title { background-color: #6699CC }
.su-spoiler.my-custom-spoiler .su-spoiler-title .su-spoiler-icon,
.su-spoiler.su-spoiler-closed.my-custom-spoiler .su-spoiler-title .su-spoiler-icon {
left: 3px;
background-color: #fff;
}
.su-spoiler.my-custom-spoiler .su-spoiler-content { background-color: #eeeeee }
.su-spoiler-title {color: #000000}
#box2
{
    height: 40px;
    width: 580px;
    background: #073763;
    font-size: 18px;
    font-style: "Roboto", sans-serif;
    color: #FFF;
    text-align: center;
    margin-top: 5px;
    margin-left: 5px;
    font-weight: bold;
    vertical-align: middle;
    display: table-cell;
    border-radius: 5px;
}




a:visited {
   color: grey;
}  

table.joomlatable th {
	padding: 5px 5px 5px 5px;
	background: #ebebeb;
	border-bottom: 1px solid #b4b4b4;
	font-weight : bold;
}

table.joomlatable tr.even td {
	padding: 5px 5px 5px 5px;
	background: #f0f0f0;
	border-bottom: 1px solid #dcdcdc;
}

table.joomlatable tr.odd td {
	padding: 5px 5px 5px 5px;
	background: #fafafa;
	border-bottom: 1px solid #dcdcdc;
}

.breadcrumbs span[typeof="v:Breadcrumb"]:last-child span[property="v:title"],
.breadcrumbs a[property="v:title"] {
    display: inline-block;
    padding: 0;
    margin-top: -3px;
    vertical-align: middle;    
    white-space: nowrap;
    overflow: hidden;
    text-overflow: ellipsis;
    margin-left: 0px;

}

/*
.urlaccesos {
    font-family: Roboto,sans-serif;
    background-color: none;
    font-weight: none;
    font-size: 14px;
    line-height: 1.3em;
    letter-spacing: 1px;  
    color: #000000;
    text-transform: none
} 
*/

a.one:link{
 text-decoration: none;
 font-family: Roboto,sans-serif;
 font-size: 14px;
 line-height: 1.3em;
 letter-spacing: 1px;  
 color: #000000
}
a.one:visited{
 text-decoration: none;
 font-family: Roboto,sans-serif;
 font-size: 14px;
 line-height: 1.3em;
 letter-spacing: 1px;  
 color: grey
}
/*
a.one:hover{
 text-decoration: none;
 font-family: Roboto,sans-serif;
 font-size: 14px;
 line-height: 1.3em;
 letter-spacing: 1px;  
 color: #000000
}

a.one:active{
 text-decoration: none;
 font-family: Roboto,sans-serif;
 font-size: 14px;
 line-height: 1.3em;
 letter-spacing: 1px;  
 color: #000000
}
*/



div.download10, span.download {
    background: #F5FAEB url("/wp-content/uploads/2015/06/download.png") no-repeat scroll 3px 5px;
    border-top: 1px dotted #78BE5A;
    border-bottom: 1px dotted #78BE5A;
}

div.tip10, span.tip {
    background: #FFFDEB url("/wp-content/uploads/2015/06/foco.png") no-repeat scroll 3px 5px;
    border-top: 1px dotted #FFC864;
    border-bottom: 1px dotted #FFC864;
}


div.download, span.download {
    background: #F5FAEB url("/wp-content/uploads/2015/06/download.png") no-repeat scroll 3px 5px;
    border-top: 1px dotted #78BE5A;
    border-bottom: 1px dotted #78BE5A;
}

div.tip, span.tip {
    background: #FFFDEB url("/wp-content/uploads/2015/06/foco.png") no-repeat scroll 3px 5px;
    border-top: 1px dotted #FFC864;
    border-bottom: 1px dotted #FFC864;
}	</style>
			<style type="text/css" id="wp-custom-css">
			/*
Puedes añadir tu propio CSS aquí.

Haz clic en el icono de ayuda de arriba para averiguar más.
*/		</style>
	<style type="text/css"></style>

		<!-- HTML5 shim and Respond.js IE8 support of HTML5 elements and media queries -->
		<!--[if lt IE 9]>
			<script src="//cdnjs.cloudflare.com/ajax/libs/html5shiv/3.7/html5shiv.min.js"></script>
			<script src="//cdnjs.cloudflare.com/ajax/libs/respond.js/1.3.0/respond.min.js"></script>
		<![endif]-->
	

</head>

<meta name="theme-color" content="#5499c7">

	<body id="top" class="home page-template page-template-page_composer page-template-page_composer-php page page-id-15 custom-background tribe-no-js site-layout-boxed site-enable-post-box-effects redsv">
			<nav id="mobile-nav-wrapper" role="navigation"></nav>
			<div id="off-canvas-body-inner">

				<!-- Top Bar -->

				<div id="top-bar" class="top-bar">
					<div class="container">
						<div class="row">
							<div class="col-sm-12">
								<div class="top-bar-right">

									
									<a class="site-social-icon" href="http://www.facebook.com/salud.sv" title="Síguenos en Facebook!" target="new"><i class="icon-social-facebook"></i></a><a class="site-social-icon" href="https://www.flickr.com/photos/minsal_sv/albums" title="Flickr" target="new"><i class="icon-social-flickr"></i></a><a class="site-social-icon" href="http://twitter.com/minsalud" title="Últimas noticias en Twitter!" target="new"><i class="icon-social-twitter"></i></a><a class="site-social-icon" href="http://www.youtube.com/comunicacionesminsal" title="Síguenos en Youtube!" target="new"><i class="icon-social-youtube"></i></a>
									<a class="instant-search-icon" href="#menu1"><i class="icon-entypo-search"></i></a>

<a href="http://publica.gobiernoabierto.gob.sv/institutions/ministerio-de-salud" title="Consultar Información Pública del Ministerio de Salud" target="_blank"><img src="/wp-content/uploads/2016/11/portal-transparencia.png" alt="Consultar Información Pública del Ministerio de Salud"></a>

								</div>

<div class="top-bar-right">
<div id="flags" class="size18"><ul id="sortable" class="ui-sortable" style="float:left"></ul></div><div id="google_language_translator"></div></div>



<div class="top-bar-right">

	<div class="zeno_font_resizer_container">
		<p class="zeno_font_resizer" style="text-align: center; font-weight: bold;">
			<span>
				<a href="#" class="zeno_font_resizer_minus" title="Decrease font size" style="font-size: 0.7em;">A</a>
				<a href="#" class="zeno_font_resizer_reset" title="Reset font size">A</a>
				<a href="#" class="zeno_font_resizer_add" title="Increase font size" style="font-size: 1.2em;">A</a>
			</span>
			<input type="hidden" id="zeno_font_resizer_value" value="body" />
			<input type="hidden" id="zeno_font_resizer_ownid" value="" />
			<input type="hidden" id="zeno_font_resizer_ownelement" value="" />
			<input type="hidden" id="zeno_font_resizer_resizeMax" value="24" />
			<input type="hidden" id="zeno_font_resizer_resizeMin" value="10" />
			<input type="hidden" id="zeno_font_resizer_resizeSteps" value="1.6" />
			<input type="hidden" id="zeno_font_resizer_cookieTime" value="31" />
		</p>
	</div>
	</div>

								<a id="open-mobile-nav" href="#mobile-nav" title="Buscar"><i class="icon-entypo-menu"></i></a>
								
								<nav id="top-nav-wrapper">
								<ul id="menu-superior" class="top-nav list-unstyled clearfix"><li id="nav-menu-item-4" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom current-menu-item current_page_item menu-item-home"><a href="http://www.salud.gob.sv/" class="menu-link main-menu-link"><span>INICIO</span></a></li>
<li id="nav-menu-item-426" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="https://mail.salud.gob.sv" class="menu-link main-menu-link"><span>CORREO</span></a></li>
<li id="nav-menu-item-3109" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/" class="menu-link main-menu-link"><span>Noticias</span></a></li>
<li id="nav-menu-item-2556" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>UACI</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-22126" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/adquisiciones-y-contrataciones-2018/" class="menu-link sub-menu-link"><span>Año 2018</span></a></li>
	<li id="nav-menu-item-14272" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/adquisiciones-y-contrataciones-2017/" class="menu-link sub-menu-link"><span>Año 2017</span></a></li>
	<li id="nav-menu-item-5653" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/adquisiciones-y-contrataciones-2016/" class="menu-link sub-menu-link"><span>Año 2016</span></a></li>
	<li id="nav-menu-item-5654" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-adquisiciones-y-contrataciones-institucional-uaci-2015/" class="menu-link sub-menu-link"><span>Año 2015</span></a></li>
	<li id="nav-menu-item-7535" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-adquisiciones-y-contrataciones-institucional-uaci-2014/" class="menu-link sub-menu-link"><span>Año 2014</span></a></li>
</ul>
</li>
<li id="nav-menu-item-15647" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>Formularios</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-1824" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-post_type menu-item-object-page"><a title="Denuncie las violaciones a su derecho a la Salud" href="http://www.salud.gob.sv/denuncias/" class="menu-link sub-menu-link"><span>DENUNCIAS A LA SALUD</span></a></li>
	<li id="nav-menu-item-15649" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/contactenos-unidad-por-el-derecho-a-la-salud/" class="menu-link sub-menu-link"><span>Unidad por el Derecho a la Salud</span></a></li>
	<li id="nav-menu-item-15652" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/hoja-de-solicitud-centro-de-capacitaciones-multiples/" class="menu-link sub-menu-link"><span>Solicitud Centro de Capacitación Max Bloch</span></a></li>
	<li id="nav-menu-item-15650" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/webmaster/" class="menu-link sub-menu-link"><span>Webmaster</span></a></li>
</ul>
</li>
<li id="nav-menu-item-6681" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>Sitio Anterior</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-6682" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/noticias-ciudadanosas-2/" class="menu-link sub-menu-link"><span>Noticias</span></a></li>
	<li id="nav-menu-item-6691" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/documentos/" class="menu-link sub-menu-link"><span>Documentos</span></a></li>
	<li id="nav-menu-item-6695" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="http://www.salud.gob.sv/galeria-de-imagenes/" class="menu-link sub-menu-link"><span>Galería de Imagenes</span></a></li>
	<li id="nav-menu-item-6699" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/audio-2/" class="menu-link sub-menu-link"><span>Audio</span></a></li>
</ul>
</li>
</ul>								</nav>
								
							</div>
						</div>
					</div>
				</div>
				<!-- End Top Bar -->
				
				<!-- Main Bar -->
								<header class="main-bar header-layout-left-logo">
					<div class="container">
						<div class="row">
							<div class="col-sm-12">

								<div id="logo" class="">

									<a href="http://www.salud.gob.sv/">

																													<img src="http://www.salud.gob.sv/wp-content/uploads/2018/02/banner_web_wpminsal_2018_V10.png" alt="MINSAL" class="logo-original" />
																	
									</a>


								</div>


																
							</div>
						</div>

					</div>
<!--META SLIDER CARRUSEL-->
<!--
<img name="banner_web_wpminsal_tres_anios_gobierno_2017" src="/wp-content/uploads/2017/05/banner_web_wpminsal_tres_anios_gobierno_2017.png" width="1200" height="170" border="0" id="banner_web_wpminsal_tres_anios_gobierno_2017" usemap="#m_banner_web_wpminsal_tres_anios_gobierno_2017" alt="" /><map name="m_banner_web_wpminsal_tres_anios_gobierno_2017" id="m_banner_web_wpminsal_tres_anios_gobierno_2017">
<area shape="rect" coords="857,0,1199,170" href="http://www.presidencia.gob.sv" target="_blank" title="www.presidencia.gob.sv" alt="www.presidencia.gob.sv" />
<area shape="rect" coords="0,0,857,170" href="http://www.salud.gob.sv" target="_parent" title="Sitio Web Ministerio de Salud de El Salvador" alt="Sitio Web Ministerio de Salud de El Salvador" />
</map>
-->

<!--
<a href="http://www.salud.gob.sv" title="Web MINSAL El Salvador" alt="Web MINSAL El Salvador">
<img src="/wp-content/uploads/2016/11/banner_web_wpminsal_2016V8.png" width="1200" height="170" border="0"></a>
-->

<!--FIN META SLIDER CARRUSEL-->

				</header>
				<!-- End Main Bar -->
				<!-- Main Navigation Bar -->
				<div class="main-nav-bar header-layout-left-logo">
					<div class="container">
						<div class="row">
							<div class="col-sm-12">
								<nav id="main-nav-wrapper"><ul id="menu-principal" class="main-nav list-unstyled"><li id="nav-menu-item-6" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>INSTITUCION</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-4299" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/estructura-organizativa/" class="menu-link sub-menu-link"><span>Estructura Organizativa</span></a></li>
	<li id="nav-menu-item-4035" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/category/institucion/area-interna/" class="menu-link sub-menu-link"><span>Área Interna</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-1033" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="https://mail.salud.gob.sv/" class="menu-link sub-menu-link"><span>Correo Institucional</span></a></li>
		<li id="nav-menu-item-2184" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/directorio-telefonico/" class="menu-link sub-menu-link"><span>Directorio Telefónico</span></a></li>
		<li id="nav-menu-item-2223" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://asp.salud.gob.sv/regulacion/default.asp" class="menu-link sub-menu-link"><span>Centro Virtual de Documentación</span></a></li>
		<li id="nav-menu-item-2227" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/biblioteca-virtual-desastres/" class="menu-link sub-menu-link"><span>Biblioteca Virtual Desastres</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-4036" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/category/institucion/marco-institucional/" class="menu-link sub-menu-link"><span>Marco Institucional</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-2190" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/historia/" class="menu-link sub-menu-link"><span>Historia</span></a></li>
		<li id="nav-menu-item-2195" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/filosofia/" class="menu-link sub-menu-link"><span>Filosofía</span></a></li>
		<li id="nav-menu-item-2232" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/autoridades/" class="menu-link sub-menu-link"><span>Autoridades</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-2256" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/otras-instituciones/" class="menu-link sub-menu-link"><span>Otras Instituciones</span></a></li>
</ul>
</li>
<li id="nav-menu-item-7" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>SERVICIOS</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-4037" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/guia/" class="menu-link sub-menu-link"><span>Guía</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-2416" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://www.salud.gob.sv/category/servicios/guia/ciudadanoa/" class="menu-link sub-menu-link"><span>Ciudadano/a</span></a></li>
		<li id="nav-menu-item-2541" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/empresas/" class="menu-link sub-menu-link"><span>Empresas</span></a></li>
		<li id="nav-menu-item-2563" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/funcionarioa/" class="menu-link sub-menu-link"><span>Funcionario/a</span></a></li>
		<li id="nav-menu-item-2612" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/ofertas-de-empleo/" class="menu-link sub-menu-link"><span>Ofertas de Empleo</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-4038" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/en-linea/" class="menu-link sub-menu-link"><span>En Línea</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-23877" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://asp.salud.gob.sv/regulacion/default.asp" class="menu-link sub-menu-link"><span>Centro Virtual de Documentación Regulatoria</span></a></li>
		<li id="nav-menu-item-2267" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa" class="menu-link sub-menu-link"><span>Guía de Servicios</span></a></li>
		<li id="nav-menu-item-2270" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/sistemas-en-linea/" class="menu-link sub-menu-link"><span>Sistemas en Línea</span></a></li>
		<li id="nav-menu-item-2273" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://saber.salud.gob.sv/" class="menu-link sub-menu-link"><span>Aula Virtual</span></a></li>
		<li id="nav-menu-item-2276" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://bbb.salud.gob.sv/" class="menu-link sub-menu-link"><span>Plataforma Webconferencia</span></a></li>
		<li id="nav-menu-item-1416" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://www.salud.gob.sv/category/servicios/en-linea/teleconferencias/" class="menu-link sub-menu-link"><span>Teleconferencias</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-6465" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/multimedia/" class="menu-link sub-menu-link"><span>Multimedia</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-5777" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/audio/" class="menu-link sub-menu-link"><span>Audio</span></a></li>
		<li id="nav-menu-item-5779" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="https://www.flickr.com/photos/minsal_sv/albums" class="menu-link sub-menu-link"><span>Fotos</span></a></li>
		<li id="nav-menu-item-14092" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/category/servicios/multimedia/videos/" class="menu-link sub-menu-link"><span>Videos</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-5974" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/documentos-institucionales/" class="menu-link sub-menu-link"><span>Documentos Institucionales</span></a></li>
</ul>
</li>
<li id="nav-menu-item-8" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>TEMAS</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-4039" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/servicios-de-salud/" class="menu-link sub-menu-link"><span>Servicios de Salud</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-3214" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/direccion-de-enfermedades-infecciosas/" class="menu-link sub-menu-link"><span>Dirección de Enfermedades Infecciosas</span></a></li>
		<li id="nav-menu-item-3221" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/programas-de-atencion-en-salud-integral-a-la-familia/" class="menu-link sub-menu-link"><span>Programas de Atención en Salud</span></a></li>
		<li id="nav-menu-item-3352" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://www.salud.gob.sv/category/temas/servicios-de-salud/sibasi/" class="menu-link sub-menu-link"><span>SIBASI</span></a></li>
		<li id="nav-menu-item-3230" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-enfermeria/" class="menu-link sub-menu-link"><span>Unidad de Enfermería</span></a></li>
		<li id="nav-menu-item-4912" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-cancer/" class="menu-link sub-menu-link"><span>Unidad de Cáncer</span></a></li>
		<li id="nav-menu-item-16784" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-salud-mental/" class="menu-link sub-menu-link"><span>Unidad de Salud Mental</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-4029" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/politicas-de-salud/" class="menu-link sub-menu-link"><span>Políticas de Salud</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-3494" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/direccion-de-vigilancia-sanitaria/" class="menu-link sub-menu-link"><span>Dirección de Vigilancia Sanitaria</span></a></li>
		<li id="nav-menu-item-3552" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/tecnologias-de-informacion-y-comunicaciones/" class="menu-link sub-menu-link"><span>Dirección de TICs</span></a></li>
		<li id="nav-menu-item-3592" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/direccion-de-desarrollo-de-recursos-humanos/" class="menu-link sub-menu-link"><span>Dirección de Desarrollo de RRHH</span></a></li>
		<li id="nav-menu-item-3793" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/direccion-de-regulacion-y-legislacion-en-salud/" class="menu-link sub-menu-link"><span>Dirección de Reg. y Leg. en Salud</span></a></li>
		<li id="nav-menu-item-3841" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/direccion-de-tecnologias-sanitarias-dirtecs/" class="menu-link sub-menu-link"><span>Dirección de Tecnologías Sanitarias</span></a></li>
		<li id="nav-menu-item-3854" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/promocion-de-la-salud/" class="menu-link sub-menu-link"><span>Promoción de la Salud</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-3210" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/gerencia-general-de-operaciones/" class="menu-link sub-menu-link"><span>Gerencia General de Operaciones</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-4304" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/adquisiciones-y-contrataciones/" class="menu-link sub-menu-link"><span>U. de Adquisiciones y Contrataciones</span></a></li>
		<li id="nav-menu-item-4292" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-de-abastecimientos/" class="menu-link sub-menu-link"><span>Unidad de Abastecimientos</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-3211" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/transversales/" class="menu-link sub-menu-link"><span>Transversales</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-4377" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a target="_blank" href="http://ins.salud.gob.sv/" class="menu-link sub-menu-link"><span>Instituto Nacional de Salud</span></a></li>
		<li id="nav-menu-item-4474" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-taxonomy menu-item-object-category"><a href="http://www.salud.gob.sv/category/temas/transversales/programas/" class="menu-link sub-menu-link"><span>Programas</span></a></li>
		<li id="nav-menu-item-4477" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/oficina-de-informacion-y-respuesta-oir/" class="menu-link sub-menu-link"><span>Oficina de Inf. y Resp. (OIR)</span></a></li>
		<li id="nav-menu-item-5074" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/unidad-por-el-derecho-a-la-salud/" class="menu-link sub-menu-link"><span>Unidad por el Derecho a la Salud</span></a></li>
	</ul>
</li>
	<li id="nav-menu-item-3445" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/preguntas-frecuentes/" class="menu-link sub-menu-link"><span>Preguntas Frecuentes</span></a></li>
</ul>
</li>
<li id="nav-menu-item-9" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>NOVEDADES</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-1131" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/category/convocatorias-de-prensa/" class="menu-link sub-menu-link"><span>Convocatorias de Prensa</span></a></li>
	<li id="nav-menu-item-15208" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/category/novedades/comunicados-de-prensa/" class="menu-link sub-menu-link"><span>Comunicados de Prensa</span></a></li>
	<li id="nav-menu-item-3092" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="/category/novedades/noticias/ciudadanosas/" class="menu-link sub-menu-link"><span>Noticias</span></a>
	<ul class="sub-menu menu-even sub-sub-menu menu-depth-2">
		<li id="nav-menu-item-14110" class="sub-menu-item sub-sub-menu-item menu-item-even menu-item-depth-2 menu-item menu-item-type-custom menu-item-object-custom"><a href="/noticias-ciudadanosas/" class="menu-link sub-menu-link"><span>Noticias Ciudadanos/as</span></a></li>
	</ul>
</li>
</ul>
</li>
<li id="nav-menu-item-2761" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>CONTÁCTENOS</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-2727" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/consultas/" class="menu-link sub-menu-link"><span>Consultas</span></a></li>
	<li id="nav-menu-item-2730" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/participacion-ciudadana/" class="menu-link sub-menu-link"><span>Participación Ciudadana</span></a></li>
	<li id="nav-menu-item-2733" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/cartas-de-derechos/" class="menu-link sub-menu-link"><span>Cartas de Derechos</span></a></li>
	<li id="nav-menu-item-2738" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/ubicacion/" class="menu-link sub-menu-link"><span>Ubicación</span></a></li>
	<li id="nav-menu-item-2724" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/regiones-de-salud/" class="menu-link sub-menu-link"><span>Regiones de Salud</span></a></li>
	<li id="nav-menu-item-2718" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/funcionarios/" class="menu-link sub-menu-link"><span>Funcionarios</span></a></li>
	<li id="nav-menu-item-2739" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/establecimientos/" class="menu-link sub-menu-link"><span>Establecimientos</span></a></li>
</ul>
</li>
<li id="nav-menu-item-156" class="main-menu-item  menu-item-even menu-item-depth-0 menu-item menu-item-type-custom menu-item-object-custom menu-item-has-children"><a href="#" class="menu-link main-menu-link"><span>AYUDA</span></a>
<ul class="sub-menu menu-odd  menu-depth-1">
	<li id="nav-menu-item-2815" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/ayuda-web/" class="menu-link sub-menu-link"><span>Ayuda Web</span></a></li>
	<li id="nav-menu-item-2877" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/mapa-del-sitio/" class="menu-link sub-menu-link"><span>Mapa del Sitio</span></a></li>
	<li id="nav-menu-item-2854" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/busqueda/" class="menu-link sub-menu-link"><span>Busqueda</span></a></li>
	<li id="nav-menu-item-2849" class="sub-menu-item  menu-item-odd menu-item-depth-1 menu-item menu-item-type-custom menu-item-object-custom"><a href="/politica-web/" class="menu-link sub-menu-link"><span>Política Web</span></a></li>
</ul>
</li>
</ul></nav>							</div>
						</div>
					</div>
				</div>
				<!-- End Main Navigation Bar -->

	
<div id="page-wrapper" class="container">
	<div class="row vwpc-row"><div class="vwpc-section-1_sidebars"><div class="col-sm-12"><hr class="section-hr"></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr"><div class="pf-content"><div class="row vwpc-row">
<div id="box1" class="col-sm-4">
<img src="/images/icon_formulario1.png"> <a href="denuncias/" title="Denuncie aquí las violaciones a su derecho a la Salud">Formulario Denuncias a la Salud</a>
</div>
<div id="box1" class="col-sm-4">
<img src="/images/icon_formulario1.png"> <a href="http://cnfv.salud.sv"  target="_blank" title="Farmacovigilancia - CNFV">Farmacovigilancia &#8211; CNFV</a>
</div>
<div id="box1" class="col-sm-4">
<img src="/images/icon_formulario1.png"> <a href="/archivos/pdf/Formularios/Lactancia_Materna/Formulario_del_derecho_a_lactar.pdf" target="_blank" title="Formulario del Derecho a Lactar">Formulario del Derecho a Lactar</a>
</div>
</div>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr"><div class="pf-content"><div class="row vwpc-row" style="background-color: #fcf3cf;">
<div class="col-sm-12" style="margin-top:20px; margin-left:0px; margin-right:0px; margin-bottom:5px;">
<div data-uk-slideset="{autoplay: true ,default: 1,small: 1,medium: 1,large: 3,xlarge: 3}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-3 uk-grid-width-xlarge-1-3">
        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><!--
Transmisión en Vivo Telesalud 2018
<div align="center">
<a href="https://bbb.salud.gob.sv/bbb/publico/create.jsp?action=invite&meetingID=Fiebre+Tifoidea" target="_blank" title="Transmisión en Vivo"><img src="/images/telesalud_2018/showbiz_boton_top_transmision_telesalud_en_vivo_wp.png"></a>
</div>
-->

<div align="center">
<a href="/programacion-de-teleconferencias-telesalud-2018/" title="Programacion de las Webconferencias 2018"><img src="/images/telesalud_2018/showbiz_boton_programacion_teleconferencias_telesalud_wp.png"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a href="http://www.empleospublicos.gob.sv/" target="_blank" title="Empleos Publicos El Salvador"><img src="/wp-content/uploads/2017/08/showbiz_boton_empleos_publicos_el_salvador_wp.png"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a href="/teleamigo/"><img src="/wp-content/uploads/2017/06/showbiz_boton_top_teleamigo_wp.png" title="TELEAMIGO 2591-7474"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a href="https://sisam.salud.gob.sv/admin/login?_moduleSelection=1" target="_blank" title="Módulo de Gestión y Control de Alimentos y Bebidas"><img src="/wp-content/uploads/2017/06/showbiz_boton_top_alimentos_bebidas_wp.png"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a href="/caja-de-herramientas-de-materiales-educativos/" title="Caja de Herramientas | Materiales Educativos"><img src="/wp-content/uploads/2017/06/showbiz_boton_top_caja_de_herramientas_wp.png"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a href="http://asp.salud.gob.sv/regulacion/default.asp" target="_blank" title="Centro Virtual de Documentación Regulatoria"><img src="/wp-content/uploads/2017/06/showbiz_boton_top_cvdr_wp.png"></a>
</div></div>
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
</div>
</div>
</div></div></div></div><div class="row vwpc-row">		<div class="vwpc-section-featured_post_slider  has-sidebar ">
						<div class="col-sm-7 col-md-8">
							<hr class="section-hr">
				<div class="flexslider no-control-nav post-slider">
	<ul class="slides">

			<li>
			<a href="http://www.salud.gob.sv/15-03-2018-nueva-area-de-pediatria-en-hospital-nacional-de-santa-ana-beneficia-a-350-mil-ninas-y-ninos/" title="Permalink to [ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños" rel="bookmark">
				<div class="post-thumbnail-wrapper">
					<img width="1140" height="641" src="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento15022018g-1140x641.jpg" class="attachment-vw_large size-vw_large wp-post-image" alt="" />				</div>

				<div class="post-box-inner">
					
					<h3 class="title">
						<span class="super-title">15 marzo, 2018</span>
						<span>[ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños</span>
					</h3>
					<span class="read-more label label-large">
						Leer Más <i class="icon-entypo-right-open"></i>
					</span>
				</div>
			</a>
		</li>
			<li>
			<a href="http://www.salud.gob.sv/07-03-2018-minsal-desarrolla-jornada-rinones-y-salud-de-las-mujeres/" title="Permalink to [ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”" rel="bookmark">
				<div class="post-thumbnail-wrapper">
					<img width="1140" height="641" src="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento07032018e-1140x641.jpg" class="attachment-vw_large size-vw_large wp-post-image" alt="" />				</div>

				<div class="post-box-inner">
					
					<h3 class="title">
						<span class="super-title">7 marzo, 2018</span>
						<span>[ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”</span>
					</h3>
					<span class="read-more label label-large">
						Leer Más <i class="icon-entypo-right-open"></i>
					</span>
				</div>
			</a>
		</li>
			<li>
			<a href="http://www.salud.gob.sv/27-02-2018-ministerio-de-salud-inicia-desparasitacion-en-poblacion-escolar/" title="Permalink to [ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar" rel="bookmark">
				<div class="post-thumbnail-wrapper">
					<img width="1140" height="641" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento27022018b-1140x641.jpg" class="attachment-vw_large size-vw_large wp-post-image" alt="" />				</div>

				<div class="post-box-inner">
					
					<h3 class="title">
						<span class="super-title">27 febrero, 2018</span>
						<span>[ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar</span>
					</h3>
					<span class="read-more label label-large">
						Leer Más <i class="icon-entypo-right-open"></i>
					</span>
				</div>
			</a>
		</li>
			<li>
			<a href="http://www.salud.gob.sv/26-02-2018-candidatas-de-santa-ana-firman-declaratoria-mas-mujeres-mas-igualdad/" title="Permalink to [ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad" rel="bookmark">
				<div class="post-thumbnail-wrapper">
					<img width="1140" height="641" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento26022018f-1140x641.jpg" class="attachment-vw_large size-vw_large wp-post-image" alt="" />				</div>

				<div class="post-box-inner">
					
					<h3 class="title">
						<span class="super-title">26 febrero, 2018</span>
						<span>[ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad</span>
					</h3>
					<span class="read-more label label-large">
						Leer Más <i class="icon-entypo-right-open"></i>
					</span>
				</div>
			</a>
		</li>
			<li>
			<a href="http://www.salud.gob.sv/22-02-2018-minsal-lanza-modelo-de-atencion-para-la-persona-adulta-mayor/" title="Permalink to [ 22-02-2018 ] MINSAL lanza modelo de atención para la persona adulta mayor" rel="bookmark">
				<div class="post-thumbnail-wrapper">
					<img width="1140" height="641" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento22022018-1140x641.jpg" class="attachment-vw_large size-vw_large wp-post-image" alt="" />				</div>

				<div class="post-box-inner">
					
					<h3 class="title">
						<span class="super-title">22 febrero, 2018</span>
						<span>[ 22-02-2018 ] MINSAL lanza modelo de atención para la persona adulta mayor</span>
					</h3>
					<span class="read-more label label-large">
						Leer Más <i class="icon-entypo-right-open"></i>
					</span>
				</div>
			</a>
		</li>
		
	</ul>
</div>			
								<div class="vwpc-section-featured_post_slider-headline row">
											<div class="post-box-wrapper col-sm-6 col-md-4 "><article class="post-24096 post-box post-box-headline">

	<h3 class="title title-small"><a href="http://www.salud.gob.sv/21-02-2018-directora-del-banco-mundial-para-centroamerica-visita-centro-nacional-de-radioterapia/" title="Permalink to [ 21-02-2018 ] Directora del Banco Mundial para Centroamérica visita Centro Nacional de Radioterapia" rel="bookmark">[ 21-02-2018 ] Directora del Banco Mundial para Centroamérica visita Centro Nacional de Radioterapia</a></h3>
	<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
		<a href="http://www.salud.gob.sv/21-02-2018-directora-del-banco-mundial-para-centroamerica-visita-centro-nacional-de-radioterapia/" class="post-date" title="Permalink to [ 21-02-2018 ] Directora del Banco Mundial para Centroamérica visita Centro Nacional de Radioterapia" rel="bookmark">21 febrero, 2018</a>
	</div>
			<div class="post-thumbnail-wrapper vw-imgliquid">
			<a href="http://www.salud.gob.sv/21-02-2018-directora-del-banco-mundial-para-centroamerica-visita-centro-nacional-de-radioterapia/" title="Permalink to [ 21-02-2018 ] Directora del Banco Mundial para Centroamérica visita Centro Nacional de Radioterapia" rel="bookmark">
				<img width="360" height="200" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento21022018e-360x200.jpg" class="attachment-vw_small size-vw_small wp-post-image" alt="" />			</a>
		</div>
	
</article></div>
											<div class="post-box-wrapper col-sm-6 col-md-4 "><article class="post-24127 post-box post-box-headline">

	<h3 class="title title-small"><a href="http://www.salud.gob.sv/14-02-2018-finaliza-segundo-curso-de-cuidados-paliativos/" title="Permalink to [ 14-02-2018 ] Finaliza Segundo “Curso de Cuidados Paliativos”" rel="bookmark">[ 14-02-2018 ] Finaliza Segundo “Curso de Cuidados Paliativos”</a></h3>
	<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
		<a href="http://www.salud.gob.sv/14-02-2018-finaliza-segundo-curso-de-cuidados-paliativos/" class="post-date" title="Permalink to [ 14-02-2018 ] Finaliza Segundo “Curso de Cuidados Paliativos”" rel="bookmark">14 febrero, 2018</a>
	</div>
			<div class="post-thumbnail-wrapper vw-imgliquid">
			<a href="http://www.salud.gob.sv/14-02-2018-finaliza-segundo-curso-de-cuidados-paliativos/" title="Permalink to [ 14-02-2018 ] Finaliza Segundo “Curso de Cuidados Paliativos”" rel="bookmark">
				<img width="360" height="200" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento14022018g-360x200.jpg" class="attachment-vw_small size-vw_small wp-post-image" alt="" />			</a>
		</div>
	
</article></div>
											<div class="post-box-wrapper col-sm-6 col-md-4 hidden-sm"><article class="post-23863 post-box post-box-headline">

	<h3 class="title title-small"><a href="http://www.salud.gob.sv/12-02-2018-minsal-recomienda-aplicar-medidas-higienicas-para-evitar-fiebre-tifoidea/" title="Permalink to [ 12-02-2018 ] MINSAL recomienda aplicar medidas higiénicas para evitar fiebre tifoidea" rel="bookmark">[ 12-02-2018 ] MINSAL recomienda aplicar medidas higiénicas para evitar fiebre tifoidea</a></h3>
	<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
		<a href="http://www.salud.gob.sv/12-02-2018-minsal-recomienda-aplicar-medidas-higienicas-para-evitar-fiebre-tifoidea/" class="post-date" title="Permalink to [ 12-02-2018 ] MINSAL recomienda aplicar medidas higiénicas para evitar fiebre tifoidea" rel="bookmark">12 febrero, 2018</a>
	</div>
			<div class="post-thumbnail-wrapper vw-imgliquid">
			<a href="http://www.salud.gob.sv/12-02-2018-minsal-recomienda-aplicar-medidas-higienicas-para-evitar-fiebre-tifoidea/" title="Permalink to [ 12-02-2018 ] MINSAL recomienda aplicar medidas higiénicas para evitar fiebre tifoidea" rel="bookmark">
				<img width="360" height="200" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento12022018_tifoidea-360x200.jpg" class="attachment-vw_small size-vw_small wp-post-image" alt="" />			</a>
		</div>
	
</article></div>
										</div>

							</div>
						<div class="col-sm-5 col-md-4">
				<aside class="sidebar-wrapper">
					<div class="sidebar-inner">
						<hr class="section-hr">
						<div id="custom_html-4" class="widget_text widget vw-sidebar-page widget_custom_html"><h3 class="widget-title">Avisos Importantes</h3><div class="textwidget custom-html-widget"><hr>

<div data-uk-slideset="{duration: 600,autoplay: true ,autoplayInterval: 10000,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://asp.salud.gob.sv/regulacion/pdf/docpublicos/Politica_Nacional_de_Salud_Mental_032018.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/banner_politica_nacional_de_salud_mental_consulta_publica-3433141905.png" alt="Banner Política Nacional de Salud Mental Consulta Pública" width="369" height="167"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://ins.salud.gob.sv/wp-content/uploads/2018/01/Bases_2018_PNM.pdf" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2018/01/banner_Premio_Nacional_de_Medicina_2018.png" title="Convocatoria 2018 | Premio Nacional de Medicina &quot;Dr. Luis Edmundo Vásquez&quot;" alt="Convocatoria 2018 | Premio Nacional de Medicina &quot;Dr. Luis Edmundo Vásquez&quot;" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://ins.salud.gob.sv/wp-content/uploads/2018/01/Gui%CC%81a_bases_PNM_2018.pdf" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2018/02/banner_Guia_Bases_PNM_2018.png" title="Guía para presentación de trabajos cientificos Premio Nacional de Medicina 2018 &quot;Dr. Luis Edmundo Vásquez&quot;" alt="Guía para presentación de trabajos cientificos Premio Nacional de Medicina 2018 &quot;Dr. Luis Edmundo Vásquez&quot;" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://ins.salud.gob.sv/wp-content/uploads/2018/01/Convocatoria_PNO.pdf" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2018/02/banner_Premio_Nacional_de_Odontologia_2018.png" title="Convocatoria 2018 | Certamen Anual de Investigación Odontológica &quot;Dr. José Benjamín Zavaleta&quot;" alt="Convocatoria 2018 |  Certamen Anual de Investigación Odontológica &quot;Dr. José Benjamín Zavaleta&quot;" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://ins.salud.gob.sv/wp-content/uploads/2018/01/Gui%CC%81a.pdf" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2018/02/banner_Guia_Bases_PNO_2018.png" title="Guía para presentación de trabajos cientificos Certamen anual de investigación odontológica 2018 &quot;Dr. José Benjamín Zavaleta&quot;" alt="Guía para presentación de trabajos cientificos Certamen anual de investigación odontológica 2018 &quot;Dr. José Benjamín Zavaleta&quot;" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://www.isss.gob.sv/index.php?option=com_content&view=article&id=1608%25regimen-especial-para-salvadorenos-en-el-exterior&catid=103%25noticias-ciudadano&Itemid=77" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2017/12/Banner_ISSS_Regimen_Salud_503_avisos_carrusel.png" title="ISSS | Régimen Salud 503" alt="ISSS | Régimen Salud 503" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/wp-content/uploads/2017/06/afiche_desinfeccion_agua_frutas_y_verduras_con_puriagua_791x1024_v062017.jpg" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/banner_desinfeccion_de_agua_frutas_y_verduras_v2_062017-beae12d51a.png" alt="Banner Desinfección de Agua Frutas y Verduras 2017" width="369" height="167"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><div align="center">
<a data-rokbox="" href="/archivos/pdf/promocion_salud/material_educativo/afiches_higiene/afiche_higiene_es_la_clave.png" data-rokbox="transitionIn:elastic;transitionOut:elastic"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2017/05/banner_higiena_es_la_clave.png" alt="Banner MINSAL Emergencias Medidas Higienicas" border="0" /></a>
</div></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="/concursos-externos/"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2016/07/banner_concursos_externos.png" title="Concursos EXternos | MINSAL" alt="Concursos Externos | MINSAL" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="/dengue/"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2016/02/banner_dengue_chiv_zika_2016wp.png" title="Campaña Dengue, Chikungunya y Zika" alt="Campaña Dengue, Chikungunya y Zika" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/promocion_salud/folleto-cuidemos-el-agua-y-eliminemos-criaderos-zancudos.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/banner_folleto_orientador_manejo_agua_reproduccion_zacudo-d33f4fb437.png" alt="Banner Folleto Orientador Manejo Agua Reproduccion Zacudo" width="369" height="167"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="/caja-de-herramientas-de-materiales-educativos/"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2016/08/banner-caja-de-herramientas.jpg" title="Caja de Herramientas de Materiales Educativos" alt="" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="/wp-content/uploads/2017/09/Comunicado-del-ISSS-Sector-Publico-Seccion-subsidios.pdf" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2017/09/banner_aviso_importante_ISSS_seccion_subsidios.png" title="AVISO IMPORTANTE | SECTOR PUBLICO - ISSS SECCION SUBSIDIOS"  alt="AVISO IMPORTANTE | SECTOR PUBLICO - ISSS SECCION SUBSIDIOS" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="https://docs.google.com/document/d/13XoHX0YEq7BTht0uTotDUFdnxHQboiOsZeOJCEj4huA/edit?usp=sharing" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2017/10/banner_catalogo_equipos_computacion_y_afines.png" title="Catálogo de equipos de computación y afines" alt="Catálogo de equipos de computación y afines" border="0" /></a></div>
                    
                    
                    
                </div>

            </li>

                </ul>

        
    </div>

    
        <ul class="uk-slideset-nav uk-dotnav uk-flex-center uk-margin-bottom-remove"></ul>
    
    
</div>

<hr></div></div><div id="custom_html-5" class="widget_text widget vw-sidebar-page widget_custom_html"><h3 class="widget-title">Accesos Directos</h3><div class="textwidget custom-html-widget"><hr>

<table id="tablepress-5" class="tablepress tablepress-id-5">
<tbody class="row-hover">
<tr class="row-1 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_siis.png"></div></td><td class="column-2"><a href="http://asp.salud.gob.sv/regulacion/default.asp" target="_blank" title="Centro Virtual de Documentación Regulatoria">Centro Virtual de Documentación</a></td>
</tr>
<tr class="row-2 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_com.png" width="21" height="19"></div></td><td class="column-2"><a href="/noticias-ciudadanosas/" title="Unidad de Comunicaciones - Noticias">Unidad de Comunicaciones - Noticias</a></td>
</tr>
<tr class="row-3 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_vig.png" width="14" height="19"></div></td><td class="column-2"><a href="/vigilancia-epidemiologica-ano-2018/" title="Vigilancia Epidemiológica 2018">Vigilancia Epidemiológica 2018</a></td>
</tr>
<tr class="row-4 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_adq.png" width="15" height="20"></div></td><td class="column-2"><a href="/boletines-epidemiologicos-2018/" title="Boletines Epidemiológicos 2018">Boletines Epidemiológicos 2018</a></td>
</tr>
<tr class="row-5 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_serv.png" width="20" height="19"></div></td><td class="column-2"><a href="/adquisiciones-y-contrataciones-2018" title="Adquisiciones y Contrataciones 2018">Adquisiciones y Contrataciones 2018</a></td>
</tr>
<tr class="row-6 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_com.png" width="21" height="19"></div></td><td class="column-2"><a href="/ofertas-de-empleo/" title="Ofertas de Empleo">Ofertas de Empleo</a></td>
</tr>
<tr class="row-7 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_siis.png"></div></td><td class="column-2"><a href="/sistemas-en-linea/" title="Sistemas en Línea">Sistemas en Línea</a></td>
</tr>
<tr class="row-8 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_saber.png"></div></td><td class="column-2"><a href="http://saber.salud.gob.sv" target="_blank" title="Centro de Conocimientos">Aula Virtual</a></td>
</tr>
<tr class="row-9 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_vac.png"></div></td><td class="column-2"><a href="/esquema-nacional-de-vacunacion-el-salvador-2017/" title="Esquema Nacional de Vacunación El Salvador 2017">Esquema Nacional de Vacunación 2017</a></td>
</tr>
<tr class="row-10 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_adq.png" width="15" height="20"></div></td><td class="column-2"><a href="/programacion-de-teleconferencias-telesalud-2018/" title="Programación de Teleconferencias 2018">Programación de Teleconferencias 2018</a></td>
</tr>
<tr class="row-11 odd">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_siis.png"></div></td><td class="column-2"><a href="/becas-cursos-congresos-diplomados-seminarios-posgrados-talleres-doctorados-maestrias-y-pasantias/" title="Becas y Cursos, Congresos, Diplomados, Seminarios, Posgrados, Talleres, Doctorados, Maestrías y Pasantías ">Becas y Cursos</a></td>
</tr>
<tr class="row-12 even">
	<td class="column-1"><div align="center"><img src="/images/slices_uno/ico_serv.png" width="20" height="19"></div></td><td class="column-2"><a href="http://rrhh.salud.gob.sv/" target="_blank" title="Observatorio de Recursos Humanos en Salud de El Salvador ">Observatorio de RRHH en Salud de El Salvador</a></td>
</tr>
</tbody>
</table>
<!-- #tablepress-5 from cache --></div></div>					</div>
				</aside>
			</div>
					</div>
		</div><div class="row vwpc-row"><div class="vwpc-section-1_sidebars"><div class="col-sm-12"><hr class="section-hr"></div></div></div><div class="row vwpc-row"><div class="vwpc-section-3_sidebars"><div class="col-sm-4"><div id="vw_widget_latest_category-10" class="widget vw-sidebar-custom-SideBarAvisos widget_vw_widget_latest_category"><h3 class="widget-title">Convocatorias de Prensa</h3><div class="post-box-list"><article class="post-24427 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/15-03-2018-0930-a-m-presidente-de-la-republica-inaugura-pabellon-de-pediatria-del-hospital-nacional-san-juan-de-dios-de-santa-ana/" title="Permalink to [15-03-2018 | 09:30 A.M.] PRESIDENTE DE LA REPÚBLICA INAUGURA PABELLÓN DE PEDIATRÍA DEL HOSPITAL NACIONAL SAN JUAN DE DIOS DE SANTA ANA" rel="bookmark">[15-03-2018 | 09:30 A.M.] PRESIDENTE DE LA REPÚBLICA INAUGURA PABELLÓN DE PEDIATRÍA DEL HOSPITAL NACIONAL SAN JUAN DE DIOS DE SANTA ANA</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/15-03-2018-0930-a-m-presidente-de-la-republica-inaugura-pabellon-de-pediatria-del-hospital-nacional-san-juan-de-dios-de-santa-ana/" class="post-date" title="Permalink to [15-03-2018 | 09:30 A.M.] PRESIDENTE DE LA REPÚBLICA INAUGURA PABELLÓN DE PEDIATRÍA DEL HOSPITAL NACIONAL SAN JUAN DE DIOS DE SANTA ANA" rel="bookmark">14 marzo, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/" title="View all posts in Convocatorias de Prensa" rel="category">Convocatorias de Prensa</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/marzo-2018/" title="View all posts in Marzo 2018" rel="category">Marzo 2018</a>		</div>
		
</article><article class="post-24281 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/07-03-2018-0830-a-m-foro-mujer-y-salud-renal/" title="Permalink to [07-03-2018 | 08:30 A.M.] FORO &#8220;MUJER Y SALUD RENAL&#8221;" rel="bookmark">[07-03-2018 | 08:30 A.M.] FORO &#8220;MUJER Y SALUD RENAL&#8221;</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/07-03-2018-0830-a-m-foro-mujer-y-salud-renal/" class="post-date" title="Permalink to [07-03-2018 | 08:30 A.M.] FORO &#8220;MUJER Y SALUD RENAL&#8221;" rel="bookmark">6 marzo, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/" title="View all posts in Convocatorias de Prensa" rel="category">Convocatorias de Prensa</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/marzo-2018/" title="View all posts in Marzo 2018" rel="category">Marzo 2018</a>		</div>
		
</article><article class="post-24166 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/27-02-2018-0900-a-m-campana-de-desparasitacion-en-poblacion-escolar/" title="Permalink to [27-02-2018 | 09:00 A.M.] CAMPAÑA DE DESPARASITACIÓN EN POBLACIÓN ESCOLAR" rel="bookmark">[27-02-2018 | 09:00 A.M.] CAMPAÑA DE DESPARASITACIÓN EN POBLACIÓN ESCOLAR</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/27-02-2018-0900-a-m-campana-de-desparasitacion-en-poblacion-escolar/" class="post-date" title="Permalink to [27-02-2018 | 09:00 A.M.] CAMPAÑA DE DESPARASITACIÓN EN POBLACIÓN ESCOLAR" rel="bookmark">26 febrero, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/" title="View all posts in Convocatorias de Prensa" rel="category">Convocatorias de Prensa</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/febrero-2018/" title="View all posts in Febrero 2018" rel="category">Febrero 2018</a>		</div>
		
</article><article class="post-24154 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/26-02-2018-1000-a-m-mujeres-santanecas-se-suman-a-declaratoria-mas-mujeres-mas-igualdad/" title="Permalink to [26-02-2018 | 10:00 A.M.] MUJERES SANTANECAS SE SUMAN A DECLARATORIA: &#8220;MAS MUJERES MAS IGUALDAD&#8221;" rel="bookmark">[26-02-2018 | 10:00 A.M.] MUJERES SANTANECAS SE SUMAN A DECLARATORIA: &#8220;MAS MUJERES MAS IGUALDAD&#8221;</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/26-02-2018-1000-a-m-mujeres-santanecas-se-suman-a-declaratoria-mas-mujeres-mas-igualdad/" class="post-date" title="Permalink to [26-02-2018 | 10:00 A.M.] MUJERES SANTANECAS SE SUMAN A DECLARATORIA: &#8220;MAS MUJERES MAS IGUALDAD&#8221;" rel="bookmark">23 febrero, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/" title="View all posts in Convocatorias de Prensa" rel="category">Convocatorias de Prensa</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/convocatorias-de-prensa/febrero-2018/" title="View all posts in Febrero 2018" rel="category">Febrero 2018</a>		</div>
		
</article></div></div></div><div class="col-sm-4"><div id="custom_html-9" class="widget_text widget vw-sidebar-custom-SideBarServicios widget_custom_html"><h3 class="widget-title">Servicios</h3><div class="textwidget custom-html-widget"><div class="post-box-list" class="title title-small">
<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/archivos/pdf/alimentos/tarifa_por_servicios.pdf" title="Tarifas de pagos por servicios" target="_blank">Tarifas de pagos por servicios.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/553" title="Extensión del Certificado de libre venta" target="_blank">Extensión del Certificado de libre venta.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/554" title="Registro sanitario y/o renovación de alimentos y bebidas importadas" target="_blank">Registro sanitario y/o renovación de alimentos y bebidas importadas.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/556" title="Registro sanitario y/o renovación de alimentos y bebidas nacionales" target="_blank">Registro sanitario y/o renovación de alimentos y bebidas nacionales.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/557" title="Autorización para importar alimentos preparados, materias primas y aditivos alimentarios" target="_blank">Autorización para importar alimentos preparados, materias primas y aditivos alimentarios.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /><a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/558" title="Reconocimiento del Registro Sanitario para Miembros de la Union Aduanera" target="_blank">Reconocimiento del Registro Sanitario para Miembros de la Union Aduanera.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/559" title="Autorización de usuarios para producir o importar alcoholes" target="_blank">Autorización de usuarios para producir o importar alcoholes.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/560" title="Dictamen técnico de condiciones de manejo y almacenamiento de productos químicos" target="_blank">Dictamen técnico de condiciones de manejo y almacenamiento de productos químicos.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/561" title="Permisos de Instalación y funcionamiento Sanitario Extendido por Unidades de Salud" target="_blank">Permisos de Instalación y funcionamiento Sanitario Extendido por Unidades de Salud.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/guia-de-servicios-gaisa/672" title="Ventanilla Única de Proyectos Habitacionales" target="_blank">Ventanilla Única de Proyectos Habitacionales.</a></p>

<p><img src="http://usam.salud.gob.sv/images/ambiental/flecha.gif" border="0" width="10" height="10" align="absMiddle" /> <a class="one" href="http://usam.salud.gob.sv/index.php/servicios/en-linea/tramites-en-linea-gaisa" title="Ayuda para trámites en línea" target="_blank">Ayuda para trámites en línea.</a></p>

</div></div></div></div><div class="col-sm-4"><div id="vw_widget_latest_category-2" class="widget vw-sidebar-custom-SideBarNoticias widget_vw_widget_latest_category"><h3 class="widget-title">Noticias</h3><div class="post-box-list"><article class="post-24464 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
					<div class="post-thumbnail-wrapper">
				<a href="http://www.salud.gob.sv/15-03-2018-nueva-area-de-pediatria-en-hospital-nacional-de-santa-ana-beneficia-a-350-mil-ninas-y-ninos/" title="Permalink to [ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños" rel="bookmark">
					<img width="360" height="360" src="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento15022018g-360x360.jpg" class="attachment-vw_square_small size-vw_square_small wp-post-image" alt="" srcset="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento15022018g-360x360.jpg 360w, http://www.salud.gob.sv/wp-content/uploads/2018/03/evento15022018g-150x150.jpg 150w, http://www.salud.gob.sv/wp-content/uploads/2018/03/evento15022018g-750x750.jpg 750w" sizes="(max-width: 360px) 100vw, 360px" />				</a>
			</div>
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/15-03-2018-nueva-area-de-pediatria-en-hospital-nacional-de-santa-ana-beneficia-a-350-mil-ninas-y-ninos/" title="Permalink to [ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños" rel="bookmark">[ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/15-03-2018-nueva-area-de-pediatria-en-hospital-nacional-de-santa-ana-beneficia-a-350-mil-ninas-y-ninos/" class="post-date" title="Permalink to [ 15-03-2018 ] Nueva área de pediatría en Hospital Nacional de Santa Ana beneficia a 350 mil niñas y niños" rel="bookmark">15 marzo, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/ano-2018/marzo-2018-ano-2018/" title="View all posts in Marzo 2018" rel="category">Marzo 2018</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/" title="View all posts in Noticias Ciudadanos/as" rel="category">Noticias Ciudadanos/as</a>		</div>
		
</article><article class="post-24380 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
					<div class="post-thumbnail-wrapper">
				<a href="http://www.salud.gob.sv/07-03-2018-minsal-desarrolla-jornada-rinones-y-salud-de-las-mujeres/" title="Permalink to [ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”" rel="bookmark">
					<img width="360" height="360" src="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento07032018e-360x360.jpg" class="attachment-vw_square_small size-vw_square_small wp-post-image" alt="" srcset="http://www.salud.gob.sv/wp-content/uploads/2018/03/evento07032018e-360x360.jpg 360w, http://www.salud.gob.sv/wp-content/uploads/2018/03/evento07032018e-150x150.jpg 150w, http://www.salud.gob.sv/wp-content/uploads/2018/03/evento07032018e-750x750.jpg 750w" sizes="(max-width: 360px) 100vw, 360px" />				</a>
			</div>
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/07-03-2018-minsal-desarrolla-jornada-rinones-y-salud-de-las-mujeres/" title="Permalink to [ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”" rel="bookmark">[ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/07-03-2018-minsal-desarrolla-jornada-rinones-y-salud-de-las-mujeres/" class="post-date" title="Permalink to [ 07-03-2018 ] MINSAL desarrolla jornada “Riñones  y Salud de las Mujeres”" rel="bookmark">7 marzo, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/ano-2018/marzo-2018-ano-2018/" title="View all posts in Marzo 2018" rel="category">Marzo 2018</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/" title="View all posts in Noticias Ciudadanos/as" rel="category">Noticias Ciudadanos/as</a>		</div>
		
</article><article class="post-24227 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
					<div class="post-thumbnail-wrapper">
				<a href="http://www.salud.gob.sv/27-02-2018-ministerio-de-salud-inicia-desparasitacion-en-poblacion-escolar/" title="Permalink to [ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar" rel="bookmark">
					<img width="360" height="360" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento27022018b-360x360.jpg" class="attachment-vw_square_small size-vw_square_small wp-post-image" alt="" srcset="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento27022018b-360x360.jpg 360w, http://www.salud.gob.sv/wp-content/uploads/2018/02/evento27022018b-150x150.jpg 150w, http://www.salud.gob.sv/wp-content/uploads/2018/02/evento27022018b-750x750.jpg 750w" sizes="(max-width: 360px) 100vw, 360px" />				</a>
			</div>
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/27-02-2018-ministerio-de-salud-inicia-desparasitacion-en-poblacion-escolar/" title="Permalink to [ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar" rel="bookmark">[ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/27-02-2018-ministerio-de-salud-inicia-desparasitacion-en-poblacion-escolar/" class="post-date" title="Permalink to [ 27-02-2018 ] Ministerio de Salud inicia desparasitación en población escolar" rel="bookmark">27 febrero, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/ano-2018/febrero-2018-ano-2018/" title="View all posts in Febrero 2018" rel="category">Febrero 2018</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/" title="View all posts in Noticias Ciudadanos/as" rel="category">Noticias Ciudadanos/as</a>		</div>
		
</article><article class="post-24240 post-box fly-in animated-content post-box-small-thumbnail clearfix">
	
					<div class="post-thumbnail-wrapper">
				<a href="http://www.salud.gob.sv/26-02-2018-candidatas-de-santa-ana-firman-declaratoria-mas-mujeres-mas-igualdad/" title="Permalink to [ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad" rel="bookmark">
					<img width="360" height="360" src="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento26022018f-360x360.jpg" class="attachment-vw_square_small size-vw_square_small wp-post-image" alt="" srcset="http://www.salud.gob.sv/wp-content/uploads/2018/02/evento26022018f-360x360.jpg 360w, http://www.salud.gob.sv/wp-content/uploads/2018/02/evento26022018f-150x150.jpg 150w, http://www.salud.gob.sv/wp-content/uploads/2018/02/evento26022018f-750x750.jpg 750w" sizes="(max-width: 360px) 100vw, 360px" />				</a>
			</div>
		
		<h3 class="title title-small"><a href="http://www.salud.gob.sv/26-02-2018-candidatas-de-santa-ana-firman-declaratoria-mas-mujeres-mas-igualdad/" title="Permalink to [ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad" rel="bookmark">[ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad</a></h3>
		<div class="post-meta header-font">
						<a class="author-name" href="http://www.salud.gob.sv/author/admin/" title="View all posts by MINSAL">MINSAL</a>,
			<a href="http://www.salud.gob.sv/26-02-2018-candidatas-de-santa-ana-firman-declaratoria-mas-mujeres-mas-igualdad/" class="post-date" title="Permalink to [ 26-02-2018 ] Candidatas de Santa Ana firman declaratoria: Más Mujeres, Más Igualdad" rel="bookmark">26 febrero, 2018</a>
		</div>
		
		<div class="post-categories clearfix">
			<a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/ano-2018/febrero-2018-ano-2018/" title="View all posts in Febrero 2018" rel="category">Febrero 2018</a><a class="label label-small" href="http://www.salud.gob.sv/category/novedades/noticias/ciudadanosas/" title="View all posts in Noticias Ciudadanos/as" rel="category">Noticias Ciudadanos/as</a>		</div>
		
</article></div></div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr">			<h1 class="section-title title title-large">
				Más Documentos			</h1>
					<div class="pf-content"><div class="row vwpc-row">
<div class="col-sm-4" style="margin-top:0px;" align="center">
<img src="/images/Estrategia_Nac_Intersectorial_Prevencion_Embarazo_en_Ninas_y_en_Adolescentes_2017_2027p.png" title="Estrategia Nacional Intersectorial de Prevención del Embarazo en Niñas y en Adolescentes 2017-2027" alt="Estrategia Nacional Intersectorial de Prevención del Embarazo en Niñas y en Adolescentes 2017-2027"><br />
<div class='w3eden'><!-- WPDM Link Template: Default Template -->


<div class="wpdm-link-tpl link-btn [color]" data-durl="http://www.salud.gob.sv/download/estrategia-nacional-intersectorial-de-prevencion-del-embarazo-en-ninas-y-en-adolescentes-2017-2027/?wpdmdl=23059" >
    <div class="media">
        <div class="pull-left"><img class="wpdm_icon" alt="Icon"   src="https://www.salud.gob.sv/wp-content/plugins/download-manager/assets/file-type-icons/pdf.png" /></div>
        <div class="media-body"><strong class="ptitle">Estrategia Nacional Intersectorial de Prevención del Embarazo en Niñas y en Adolescentes 2017-2027 <span class="label label-default" style="font-weight: 400;">7.03 MB</span></strong>
            <div><strong><a class='wpdm-download-link btn btn-info btn-xs' rel='nofollow' href='#' onclick="location.href='http://www.salud.gob.sv/download/estrategia-nacional-intersectorial-de-prevencion-del-embarazo-en-ninas-y-en-adolescentes-2017-2027/?wpdmdl=23059';return false;">Descargar</a></strong></div>
        </div>
    </div>
</div>
<div style="clear: both"></div>
</div></div>
<p><!--


<div class="col-sm-4" style="margin-top:0px;" align="center">
<img src="/images/Plan_Operativo_Institucional_2017.png" title="Plan Operativo Institucional | Enero - Diciembre 2017" alt="Plan Operativo Institucional | Enero - Diciembre 2017"><br />
[wpdm_package id='15533']</div>


--></p>
<div class="col-sm-4" style="margin-top:0px;" align="center">
<img src="/images/Plan_Estrategico_Institucional_en_Salud_PEI_2014-2019.png" title="Plan Estratégico 2014-2019" alt="Plan Estratégico 2014-2019"></p>
<div class='w3eden'><!-- WPDM Link Template: Default Template -->


<div class="wpdm-link-tpl link-btn [color]" data-durl="http://www.salud.gob.sv/download/plan-estrategico-2014-2019/?wpdmdl=15531" >
    <div class="media">
        <div class="pull-left"><img class="wpdm_icon" alt="Icon"   src="https://www.salud.gob.sv/wp-content/plugins/download-manager/assets/file-type-icons/pdf.png" /></div>
        <div class="media-body"><strong class="ptitle">Plan Estratégico 2014-2019 <span class="label label-default" style="font-weight: 400;">2.03 MB</span></strong>
            <div><strong><a class='wpdm-download-link btn btn-info btn-xs' rel='nofollow' href='#' onclick="location.href='http://www.salud.gob.sv/download/plan-estrategico-2014-2019/?wpdmdl=15531';return false;">Descargar</a></strong></div>
        </div>
    </div>
</div>
<div style="clear: both"></div>
</div></div>
<div class="col-sm-4" style="margin-top:0px;" align="center">
<div data-uk-slideset="{animation: 'slide-horizontal',autoplay: true ,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><div class="uk-overlay uk-overlay-hover uk-border-rounded"><img src="/wp-content/uploads/2017/07/MINSAL_Informe_de_Labores_2016_2017_portada.png" class="uk-border-rounded" alt="MINSAL Informe De Labores 2016 2017 Portada" width="256" height="329"><a class="uk-position-cover" href="/informe-de-rendicion-de-cuentas-2016-2017/"></a></div></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><div class="uk-overlay uk-overlay-hover uk-border-rounded"><img src="/wp-content/uploads/2017/07/MINSAL_Informe_de_Labores_2015-2016_portada.png" class="uk-border-rounded" alt="MINSAL Informe De Labores 2015 2016 Portada" width="256" height="329"><a class="uk-position-cover" href="/informe-de-rendicion-de-cuentas-2015-2016/"></a></div></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
<b>Informes de Labores y Rendición de Cuentas<br />Años 2016-2017 | 2015-2016</b><br />
<!--
<a href="http://www.salud.gob.sv/informe-de-rendicion-de-cuentas-2015-2016/"><img src="/archivos/pdf/Rendicion-de-Cuentas/2015-2016/Informe_de_Labores_2015-2016_portada.png" title="Informe de Labores, Suplemento, Presentación y Video 2015-2016" alt="Informe de Labores, Suplemento, Presentación y Video 2015-2016" /></a>
-->
</div>
</div>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr"><div class="pf-content"><div class="row vwpc-row" style="background-color: #666600; ">
<div class="col-sm-3" style="margin-top:20px;">
<div data-uk-slideset="{duration: 400,autoplay: true ,autoplayInterval: 4000,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://asp.salud.gob.sv/regulacion/default.asp" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/CVDRS-fa503c8518.png" alt="Centro Virtual de Documentación Regulatoria" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://www.paho.org/resscad/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/boton_izq_XXX_RESSCAD_ELS2014-3e833c0a5d.png" alt="Boton Izq XXX RESSCAD ELS2014" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://ins.salud.gob.sv/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_insv2-ab93f604b8.png" alt="Instituto Nacional de Salud" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://www.incap.org.gt/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/boton_izq_incap-90d684c1d1.png" alt="Instituto de Nutrición de Centro América y Panamá (INCAP)" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://asp.salud.gob.sv/desastres/index2.html" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/BVDESASTRES-5187c6a917.jpg" alt="Bibliotec Virtual Desastres" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://www.teg.gob.sv/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_teg-f1b5018fdd.png" alt="Tribunal de Ética Gubernamental" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
</div>
<div class="col-sm-3" style="margin-top:20px;">
<div data-uk-slideset="{duration: 400,autoplay: true ,autoplayInterval: 4000,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/?p=3608"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/uploads/2015/07/becas_cursos.png" alt="Becas Cursos" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/?p=2610"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/uploads/2015/07/ofertas_de_empleo.png" alt="Ofertas De Empleo" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/programacion-de-teleconferencias-2017/"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/uploads/2017/10/teleconferencias.png" alt="Teleconferencias2016" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                    
                    
                    
                    
                    
                                        <div class="uk-margin"><a href="http://cnfv.salud.sv/" target="_blank"><img style="display: block; margin-left: auto; margin-right: auto;" src="/wp-content/uploads/2017/10/logo_CNFV_carrusel_minsal.png" title="Farmacovigilancia -CNFV"  alt="Farmacovigilancia -CNFV" style="border: 1px solid #eee; -webkit-border-radius: 10px; -moz-border-radius: 10px; border-radius: 10px; margin-bottom:10px;"></a></div>
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/unidad-reguladora-y-asesora-de-radiaciones/"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/uploads/2015/07/logo_UNRA.jpg" alt="Logo UNRA" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
</div>
<div class="col-sm-3" style="margin-top:20px;">
<div data-uk-slideset="{duration: 400,autoplay: true ,autoplayInterval: 4000,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/politica-nacional-de-salud-2015-2019_version_imprenta.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/politica_nac_salud_2015-2019-46ec94dda4.png" alt="Politica Nac Salud 2015 2019" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://asp.salud.gob.sv/regulacion/pdf/planes/Plan_Estrategico_Institucional_en_Salud_PEI_2014-2019.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/PEI2014-2019_MINSAL_bottom-5f816fd32a.png" alt="PEI2014 2019 MINSAL Bottom" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Documentos_Externos/COMISCA-SICA/Politica-Regional-de-Salud-del-SICA-2015-2022-COMISCA.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/politica-regional-de-salud-del-sica-2015-2022-comisca-0e552f0d52.png" alt="Politica Regional De Salud Del Sica 2015 2022 Comisca" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Documentos_Externos/COMISCA-SICA/Plan-de-Salud-de-Centroamerica-y-Republica-Dominicana-2016-2020-COMISCA.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/plan-de-salud-CA-RD-2016-2020-comisca-eda7446987.png" alt="Plan De Salud CA RD 2016 2020 Comisca" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Documentos_Externos/COMISCA-SICA/Agenda-de-Salud-de-Centroamerica-y-Republica-Dominicana-2009-2018-COMISCA.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/agenda-de-salud-CA-RD-2009-2018-8ae5a1a42b.png" alt="Agenda De Salud CA RD 2009 2018" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Suplemento_La_Reforma_de_Salud_Avanza.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/carrusel_Suplemento_La_Reforma_de_Salud_Avanza_bottom-4610287f5c.png" alt="Carrusel Suplemento La Reforma De Salud Avanza Bottom" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Estudio_Nac_de_Yoduria_2012_Unidad_Nutrucion.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/portada_estudio_yoduria2012-f843395146.png" alt="Estudio Nacional de Yoduria | El Salvador, Agosto - Octubre 2012" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Encuesta_Nacional_de_Salud_ENS-2014.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/portada_ENS2014-28c31f9483.png" alt="Portada ENS2014" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="/archivos/pdf/Encuesta_mundial_salud_escolar_el_salvador2014.pdf" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/encuesta_escolar-4610287f5c.png" alt="Encuesta Escolar" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
</div>
<div class="col-sm-3" style="margin-top:20px;">
<div data-uk-slideset="{duration: 400,autoplay: true ,autoplayInterval: 4000,default: 1,small: 1,medium: 1,large: 1,xlarge: 1}">

    
    <div class="uk-slidenav-position uk-margin">

        <ul class="uk-slideset uk-grid uk-grid-match uk-flex-center uk-grid-width-1-1 uk-grid-width-small-1-1 uk-grid-width-medium-1-1 uk-grid-width-large-1-1 uk-grid-width-xlarge-1-1">
        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://publica.gobiernoabierto.gob.sv/institutions/ministerio-de-salud" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_portal_transparencia_MINSAL_carrusel-adc9579e60.png" alt="Portal de Transparencia MINSAL" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://infoutil.gobiernoabierto.gob.sv/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo-infoUtil-8067feb4d6.png" alt="Logo InfoUtil" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://elsalvador.eregulations.org/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_infotramites-a6fdf31451.png" alt="Logo Infotramites" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="https://www.miempresa.gob.sv/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_miempresa-a6fdf31451.png" alt="Logo Miempresa" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

        
            <li>

                <div class="uk-panel uk-text-center">

                                        <a class="uk-position-cover uk-position-z-index" href="http://premiocalidad.presidencia.gob.sv/" target="_blank"></a>
                    
                    
                                        <div class="uk-text-center uk-panel-teaser"><img src="/wp-content/plugins/widgetkit/cache/logo_ESCalidad-8067feb4d6.png" alt="Logo ESCalidad" width="170" height="121"></div>
                    
                    
                    
                    
                    
                    
                </div>

            </li>

                </ul>

                <a href="#" class="uk-slidenav  uk-slidenav-previous uk-hidden-touch" data-uk-slideset-item="previous"></a>
        <a href="#" class="uk-slidenav  uk-slidenav-next uk-hidden-touch" data-uk-slideset-item="next"></a>
        
    </div>

    
    
    
</div>
</div>
</div>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr">			<h1 class="section-title title title-large">
				Política Nacional de Salud 2015-2019			</h1>
					<div class="pf-content"><div class="row vwpc-row">
<div class="col-sm-4" style="margin-top:0px;" align="center"><img src="/images/Poltica_Nacional_de_Salud_2015_2019_DO.png" title="Versión Diario Oficial"><br />
<div class='w3eden'><!-- WPDM Link Template: Default Template -->


<div class="wpdm-link-tpl link-btn [color]" data-durl="http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019-diario-oficial-no-182-tomo-no-413-del-03-10-2016-acuerdo-no-1422/?wpdmdl=15112" >
    <div class="media">
        <div class="pull-left"><img class="wpdm_icon" alt="Icon"   src="https://www.salud.gob.sv/wp-content/plugins/download-manager/assets/file-type-icons/pdf.png" /></div>
        <div class="media-body"><strong class="ptitle">Política Nacional de Salud 2015-2019 | Diario Oficial No.182, Tomo No.413 del 03-10-2016. Acuerdo No.1422. <span class="label label-default" style="font-weight: 400;">188.65 KB</span></strong>
            <div><strong><a class='wpdm-download-link btn btn-info btn-xs' rel='nofollow' href='#' onclick="location.href='http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019-diario-oficial-no-182-tomo-no-413-del-03-10-2016-acuerdo-no-1422/?wpdmdl=15112';return false;">Descargar</a></strong></div>
        </div>
    </div>
</div>
<div style="clear: both"></div>
</div>
</div>
<div class="col-sm-4" style="margin-top:0px;" align="center"><img src="/images/Poltica_Nacional_de_Salud_2015_2019_version_imprenta.png" title="Versión Imprenta"><br />
<div class='w3eden'><!-- WPDM Link Template: Default Template -->


<div class="wpdm-link-tpl link-btn [color]" data-durl="http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019/?wpdmdl=15109" >
    <div class="media">
        <div class="pull-left"><img class="wpdm_icon" alt="Icon"   src="https://www.salud.gob.sv/wp-content/plugins/download-manager/assets/file-type-icons/pdf.png" /></div>
        <div class="media-body"><strong class="ptitle">Política Nacional de Salud 2015-2019 | Versión Imprenta <span class="label label-default" style="font-weight: 400;">585.41 KB</span></strong>
            <div><strong><a class='wpdm-download-link btn btn-info btn-xs' rel='nofollow' href='#' onclick="location.href='http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019/?wpdmdl=15109';return false;">Descargar</a></strong></div>
        </div>
    </div>
</div>
<div style="clear: both"></div>
</div></div>
<div class="col-sm-4" style="margin-top:0px;" align="center"><img src="/images/Poltica_Nacional_de_Salud_2015_2019_version_popular.png" title="Versión Diario Popular"><br />
<div class='w3eden'><!-- WPDM Link Template: Default Template -->


<div class="wpdm-link-tpl link-btn [color]" data-durl="http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019-version-popular/?wpdmdl=15180" >
    <div class="media">
        <div class="pull-left"><img class="wpdm_icon" alt="Icon"   src="https://www.salud.gob.sv/wp-content/plugins/download-manager/assets/file-type-icons/pdf.png" /></div>
        <div class="media-body"><strong class="ptitle">Política Nacional de Salud 2015-2019 | Versión Popular <span class="label label-default" style="font-weight: 400;">32.70 MB</span></strong>
            <div><strong><a class='wpdm-download-link btn btn-info btn-xs' rel='nofollow' href='#' onclick="location.href='http://www.salud.gob.sv/download/politica-nacional-de-salud-2015-2019-version-popular/?wpdmdl=15180';return false;">Descargar</a></strong></div>
        </div>
    </div>
</div>
<div style="clear: both"></div>
</div></div>
</div>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-1_sidebars"><div class="col-sm-12"><hr class="section-hr"></div></div></div><div class="row vwpc-row"><div class="vwpc-section-3_sidebars"><div class="col-sm-4"><div id="vw_widget_custom_text-4" class="widget vw-sidebar-custom-SideBarMultimedia2 widget_vw_widget_custom_text"><h3 class="widget-title">UDECOM MINSAL 2018</h3>			<div align="center">
<!--
<iframe width="100%" height="245" src="https://www.youtube.com/embed/_wOgOhIItDw?rel=0" frameborder="0" allowfullscreen></iframe>
-->

<!--
AÑO 2017
<iframe width="100%" height="245" src="http://www.youtube.com/embed/videoseries?list=PLfQ_63-k_c8arfLdneWLcxKtRl_yy1Yq8&hl=es_ES&rel=0" name="UDECOM2017" frameborder="0" allowfullscreen></iframe>
</div>
-->

<iframe width="100%" height="245" src="http://www.youtube.com/embed/videoseries?list=PLfQ_63-k_c8Y2Ft8-V5JD4Ct9uwUR0WlN&hl=es_ES&rel=0" name="UDECOM2017" frameborder="0" allowfullscreen></iframe>
</div>




		</div></div><div class="col-sm-4"><div id="vw_widget_custom_text-7" class="widget vw-sidebar-blog widget_vw_widget_custom_text"><h3 class="widget-title">Spot de Campañas</h3>			<div align="center">
<iframe width="100%" height="245" src="https://www.youtube.com/embed/videoseries?list=PLfQ_63-k_c8ZfscBeEv-PDctdzPp7z8HR&hl=es_ES&rel=0"  name="SPOTS2017" frameborder="0" allowfullscreen></iframe>
</div>		</div></div><div class="col-sm-4"><div id="vw_widget_custom_text-5" class="widget vw-sidebar-custom-SideBarMultimedia3 widget_vw_widget_custom_text"><h3 class="widget-title">Hablemos de VIHDA</h3>			<div align="center">
<iframe width="100%" height="245" src="http://www.youtube.com/embed/videoseries?list=PLV2iO17j3vxVcqTWY4I5WCs_mu5-o2aTu&hl=es_ES&rel=0" name="HABLEMOSVIHDA" frameborder="0" allowfullscreen></iframe>
</div>
<div align="center">
<a data-rokbox="" href="/archivos/comunicaciones/programacion_Hablemos_VIHDA_2015.jpg" target="_blank" data-lightbox="transitionIn:elastic;transitionOut:elastic"><b>Ver Horarios de Transmisión</b></a>
</div>		</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr">			<h1 class="section-title title title-large">
				Empleos Públicos en El Salvador			</h1>
					<div class="pf-content"><div class="row vwpc-row">
<div class="col-sm-8">
<a href="http://www.empleospublicos.gob.sv/" title="Empleos Públicos en El Salvador" target="_blank"><img src="/wp-content/uploads/2017/07/banner_bottom_empleos_publicos_el_salvador.png" style="border: 1px solid #ccc; -webkit-border-radius: 10px; -moz-border-radius: 10px; border-radius: 10px; margin-bottom:10px;"></a><br />
<a href="http://www.empleospublicos.gob.sv/pasos.aspx" target="_blank" title="Pasos de ¿Cómo participar en un concurso? en Empleos Públicos en El Salvador "><img src="/wp-content/uploads/2017/07/bannerPasosAbajo.png"></a>
</div>
<div class="col-sm-4">
<div><iframe src="https://www.youtube.com/embed/lbAnizGrYvM" width="320" height="240" title="Tutorial de Empleos Públicos de El Salvador" frameborder="0" allowfullscreen="allowfullscreen"></iframe></div>
</div>
</div>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr">			<h1 class="section-title title title-large">
				Audios			</h1>
					<div class="pf-content"><div class="row vwpc-row">
<div class="col-sm-6" style="margin-top:0px;">
        <font face="Arial" size="5"><b>Programas de Radio ¡Viva la Salud!</b></font><br />
        <!--[if lt IE 9]><script>document.createElement('audio');</script><![endif]-->
<div class="wp-playlist wp-audio-playlist wp-playlist-light">
		<div class="wp-playlist-current-item"></div>
		<audio controls="controls" preload="none" width="1118"></audio>
	<div class="wp-playlist-next"></div>
	<div class="wp-playlist-prev"></div>
	<noscript>
	<ol><li><a href='http://www.salud.gob.sv/wp-content/uploads/2018/03/programa383_12032018.mp3'>Programa de Radio No.383 [ 12/03/2018 ]</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2018/02/programa382_05032018.mp3'>Programa de Radio No.382 [ 05/03/2018 ]</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2018/02/programa381_26022018.mp3'>Programa de Radio No.381 [ 26/02/2018 ]</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2018/02/programa380_19022018.mp3'>Programa de Radio No.380 [ 19/02/2018 ]</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2018/02/programa379_12022018.mp3'>Programa de Radio No.379 [ 12/02/2018 ]</a></li></ol>
	</noscript>
	<script type="application/json" class="wp-playlist-script">{"type":"audio","tracklist":true,"tracknumbers":true,"images":true,"artists":false,"tracks":[{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2018\/03\/programa383_12032018.mp3","type":"audio\/mpeg","title":"Programa de Radio No.383 [ 12\/03\/2018 ]","caption":"","description":"\"Programa de Radio No.383 [ 12\/03\/2018 ]\" en \u00a1Viva la Salud! por Entrevista: Dr. Carlos Orantes, Especialista en Nefrolog\u00eda y Colaborador T\u00e9cnico de la Direcci\u00f3n de Enfermedades No Transmisibles del MINSAL para hablar sobre la salud renal. G\u00e9nero: Blues.","meta":{"artist":"Entrevista: Dr. Carlos Orantes, Especialista en Nefrolog\u00eda y Colaborador T\u00e9cnico de la Direcci\u00f3n de Enfermedades No Transmisibles del MINSAL para hablar sobre la salud renal.","album":"\u00a1Viva la Salud!","genre":"Blues","length_formatted":"46:37"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2018\/02\/programa382_05032018.mp3","type":"audio\/mpeg","title":"Programa de Radio No.382 [ 05\/03\/2018 ]","caption":"","description":"\"Programa de Radio No.382 [ 05\/03\/2018 ]\" en \u00a1Viva la Salud! por Entrevsita Yanira Argueta, Directora Ejecutiva de ISDEMU para hablar sobre el D\u00eda Internacional de la Mujer.. G\u00e9nero: Blues.","meta":{"artist":"Entrevsita Yanira Argueta, Directora Ejecutiva de ISDEMU para hablar sobre el D\u00eda Internacional de la Mujer.","album":"\u00a1Viva la Salud!","genre":"Blues","length_formatted":"52:50"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2018\/02\/programa381_26022018.mp3","type":"audio\/mpeg","title":"Programa de Radio No.381 [ 26\/02\/2018 ]","caption":"","description":"\"Programa de Radio No.381 [ 26\/02\/2018 ]\" en \u00a1Viva la Salud! por Hablaremos sobre la Campa\u00f1a de Vacunaci\u00f3n Canina y Felina.","meta":{"artist":"Hablaremos sobre la Campa\u00f1a de Vacunaci\u00f3n Canina y Felina","album":"\u00a1Viva la Salud!","length_formatted":"53:50"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2018\/02\/programa380_19022018.mp3","type":"audio\/mpeg","title":"Programa de Radio No.380 [ 19\/02\/2018 ]","caption":"","description":"\"Programa de Radio No.380 [ 19\/02\/2018 ]\" en \u00a1Viva la Salud! por Entrevista Dra. Alexandra Portillo, Coordinadora de las Enfermedades Infecciosas Desatendidas del MINSAL para hablar sobre el Parasitismo.. G\u00e9nero: Blues.","meta":{"artist":"Entrevista Dra. Alexandra Portillo, Coordinadora de las Enfermedades Infecciosas Desatendidas del MINSAL para hablar sobre el Parasitismo.","album":"\u00a1Viva la Salud!","genre":"Blues","length_formatted":"55:47"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2018\/02\/programa379_12022018.mp3","type":"audio\/mpeg","title":"Programa de Radio No.379 [ 12\/02\/2018 ]","caption":"","description":"\"Programa de Radio No.379 [ 12\/02\/2018 ]\" en \u00a1Viva la Salud! por Entrevista Dr. Alvaro Hugo Salgado Rold\u00e1n, Director del Hospital Nacional Especializado de Ni\u00f1os \"Benjam\u00edn Bloom\".. G\u00e9nero: Blues.","meta":{"artist":"Entrevista Dr. Alvaro Hugo Salgado Rold\u00e1n, Director del Hospital Nacional Especializado de Ni\u00f1os \"Benjam\u00edn Bloom\".","album":"\u00a1Viva la Salud!","genre":"Blues","length_formatted":"54:03"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}}]}</script>
</div>
	
<div align="center">
       [ <a href="/audio/#VLS"><b>Escuchar más Programas de Radio</b></a> ] [ <a href="/multimedia-audio-3/#VLS"><b>Descargar Programas de Radio</b></a> ]
	</div>
</div>
<div class="col-sm-6" style="margin-top:0px;">
        <font face="Arial" size="5"><b>Cuñas de Radio | Dale Salud a tu Vida</b></font><br />
        <div class="wp-playlist wp-audio-playlist wp-playlist-light">
		<div class="wp-playlist-current-item"></div>
		<audio controls="controls" preload="none" width="1118"></audio>
	<div class="wp-playlist-next"></div>
	<div class="wp-playlist-prev"></div>
	<noscript>
	<ol><li><a href='http://www.salud.gob.sv/wp-content/uploads/2017/04/MINSAL-Dale-salud-a-tu-vida-AZUCAR-Radio-CORREGIDO.mp3'>MINSAL - Dale salud a tu vida - AZUCAR</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2017/04/MINSAL-Dale-salud-a-tu-vida-GRASAS-Radio-CORREGIDO.mp3'>MINSAL - Dale salud a tu vida - GRASAS</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2017/04/MINSAL-Dale-salud-a-tu-vida-SAL-Radio-CORREGIDO.mp3'>MINSAL - Dale salud a tu vida - SAL</a></li><li><a href='http://www.salud.gob.sv/wp-content/uploads/2017/04/MINSAL-Dale-salud-a-tu-vida-VIÑETAS-Radio-CORREGIDO.mp3'>MINSAL - Dale salud a tu vida - VIÑETAS</a></li></ol>
	</noscript>
	<script type="application/json" class="wp-playlist-script">{"type":"audio","tracklist":true,"tracknumbers":true,"images":true,"artists":true,"tracks":[{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2017\/04\/MINSAL-Dale-salud-a-tu-vida-AZUCAR-Radio-CORREGIDO.mp3","type":"audio\/mpeg","title":"MINSAL - Dale salud a tu vida - AZUCAR","caption":"","description":"\"MINSAL - Dale salud a tu vida - AZUCAR Radio CORREGIDO\". Lanzamiento: 2017. Pista 1.","meta":{"year":"2017","length_formatted":"0:30"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2017\/04\/MINSAL-Dale-salud-a-tu-vida-GRASAS-Radio-CORREGIDO.mp3","type":"audio\/mpeg","title":"MINSAL - Dale salud a tu vida - GRASAS","caption":"","description":"\"MINSAL - Dale salud a tu vida - GRASAS Radio CORREGIDO\". Lanzamiento: 2017. Pista 1.","meta":{"year":"2017","length_formatted":"0:30"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2017\/04\/MINSAL-Dale-salud-a-tu-vida-SAL-Radio-CORREGIDO.mp3","type":"audio\/mpeg","title":"MINSAL - Dale salud a tu vida - SAL","caption":"","description":"\"MINSAL - Dale salud a tu vida - SAL Radio CORREGIDO\". Lanzamiento: 2017. Pista 1.","meta":{"year":"2017","length_formatted":"0:30"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}},{"src":"http:\/\/www.salud.gob.sv\/wp-content\/uploads\/2017\/04\/MINSAL-Dale-salud-a-tu-vida-VIN\u0303ETAS-Radio-CORREGIDO.mp3","type":"audio\/mpeg","title":"MINSAL - Dale salud a tu vida - VIN\u0303ETAS","caption":"","description":"\"MINSAL - Dale salud a tu vida - VIN\u0303ETAS Radio CORREGIDO\". Lanzamiento: 2017. Pista 1.","meta":{"year":"2017","length_formatted":"0:35"},"image":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64},"thumb":{"src":"http:\/\/www.salud.gob.sv\/wp-includes\/images\/media\/audio.png","width":48,"height":64}}]}</script>
</div>
	
<div align="center">
        [ <a href="/multimedia-audio-3/#SPOT-RADIO"><b>Descargar Cuñas de Radio</b></a> ]
        </div>
</div>
</div>
<p><!--


<div class="row vwpc-row">



<div class="col-sm-6" style="margin-top:0px;">
<font face="Arial" size="5"><b>Programas de Radio ¡Viva la Salud!</b></font><br />
[playlist artists="false" ids="18411,18263,18262,17822,17552"]</div>





<div align="center">
[ <a href="/audio/#VLS"><b>Escuchar más Programas de Radio</b></a> ]</div>


</div>






<div class="col-sm-6" style="margin-top:0px;">
<font face="Arial" size="5"><b>Cuñas de Radio | Dale Salud a tu Vida</b></font><br />
[playlist ids="17128,17129,17130,17131" style="light"]</div>





<div align="center">
[ <a href="/multimedia-audio-3/#SPOT-RADIO"><b>Descargar Cuñas de Radio</b></a> ]
</div>




</div>


--></p>
</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-1_sidebars"><div class="col-sm-12"><hr class="section-hr"><div id="showbiz-widget-2" class="widget vw-sidebar-custom-SideBarMultimedia1 widget_showbiz"><h3 class="widget-title"></h3>				
			<!-- START SHOWBIZ 1.7.2 -->	
			
						
						<style type="text/css">
				/********************************************

	STYLE SETTINGS FOR THE GREY SKIN

*********************************************/

#showbiz_1_1.showbiz-container{
	max-width:1210px;
	min-width:300px;
}

#showbiz_1_1 .showbiz-title				{
                                        margin-top:10px;
                                        text-align:center;
                                    }

#showbiz_1_1 .showbiz-title,
#showbiz_1_1 .showbiz-title a,
#showbiz_1_1 .showbiz-title a:visited,
#showbiz_1_1 .showbiz-title a:hover		{
                                            color:#555;
                                            font-family: 'Open Sans', sans-serif;
                                            font-size:14px;
                                            text-transform:uppercase;
                                            text-decoration: none;
                                            font-weight:700;
                                    }

#showbiz_1_1 .showbiz-description		{
                                        margin-top:10px;
                                        text-align:center;
                                        font-size:13px;
                                        line-height:22px;
                                        color:#777;
                                        font-family: 'Open Sans', sans-serif;
                                    }



#showbiz_1_1  .mediaholder 				{	background-color:#003366;
                                        border:1px solid #f5f5f5;
                                        border-radius:2px;-moz-border-radius:2px;-webkit-border-radius:2px;
                                        padding:7px;
                                    }

#showbiz_1_1  .hovercover				{	background:rgba(0,0,0,0.5);  }

#showbiz_1_1 li:hover .mediaholder img  {	filter: url("data:image/svg+xml;utf8,<svg xmlns=\'http://www.w3.org/2000/svg\'><filter id=\'grayscale\'><feColorMatrix type=\'matrix\' values=\'0.3333 0.3333 0.3333 0 0 0.3333 0.3333 0.3333 0 0 0.3333 0.3333 0.3333 0 0 0 0 0 1 0\'/></filter></svg>#grayscale");
                                        filter: gray; /* IE6-9 */
                                        -webkit-filter: grayscale(100%);
                                    }
/*** WHITE NAV BUTTONS ***/
#showbiz_1_1 .showbiz-navigation						{	margin-bottom:20px;}

#showbiz_1_1 .sb-navigation-left,
#showbiz_1_1 .sb-navigation-right,
#showbiz_1_1 .sb-navigation-play						{	border:1px solid #000; }

#showbiz_1_1 .showbiz-navigation i						{	color:#000;   }

#showbiz_1_1 .sb-navigation-left:hover,
#showbiz_1_1 .sb-navigation-right:hover					{	border:1px solid #000;}

#showbiz_1_1 .sb-navigation-left.notclickable:hover,
#showbiz_1_1 .sb-navigation-right.notclickable:hover	{	border:1px solid #000;}
#showbiz_1_1 .sb-navigation-left, .sb-navigation-right, .sb-navigation-play {
    border-radius: 0px;
    cursor: pointer;
    display: inline-block;
    padding: 1px 3px;
    transition: all 0.3s ease-in-out 0s;
} 
				
				.showbiz-drag-mouse {
					cursor:url(http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/css/openhand.cur), move;
				}
				.showbiz-drag-mouse.dragged {
					cursor:url(http://www.salud.gob.sv/wp-content/plugins/showbiz/showbiz-plugin/css/closedhand.cur), move;
				}
			</style>
						
			<div id="showbiz_1_1" class="showbiz-container" style="margin:0px auto;margin-top:0px;margin-bottom:0px;">
				
								
				<div class="showbiz"  data-left="#showbiz_left_1" data-right="#showbiz_right_1" data-play="#showbiz_play_1" >
					<div class="overflowholder">
					
						<ul>					<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/12/logo_503_ISSS290x155.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.isss.gob.sv/index.php?option=com_content&#038;view=article&#038;id=1608%regimen-especial-para-salvadorenos-en-el-exterior&#038;catid=103%noticias-ciudadano&#038;Itemid=77#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/12/logo_503_ISSS290x155.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.isss.gob.sv/index.php?option=com_content&#038;view=article&#038;id=1608%regimen-especial-para-salvadorenos-en-el-exterior&#038;catid=103%noticias-ciudadano&#038;Itemid=77#new_tab">ISSS | Régimen Salud 503</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/03/gobernando_con_la_gente.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.presidencia.gob.sv/gobernando-con-la-gente/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/03/gobernando_con_la_gente.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.presidencia.gob.sv/gobernando-con-la-gente/#new_tab">Gobernando con la Gente</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/03/casa-abierta.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.presidencia.gob.sv/temas/casa-abierta/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/03/casa-abierta.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.presidencia.gob.sv/temas/casa-abierta/#new_tab">Casa Abierta</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/03/logo_AvancES.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://avances.sv/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/03/logo_AvancES.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://avances.sv/#new_tab">AvancES</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/03/cronica_ciudadana.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.presidencia.gob.sv/temas/cronica-salvadorena/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/03/cronica_ciudadana.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.presidencia.gob.sv/temas/cronica-salvadorena/#new_tab">Crónica Ciudadana</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2017/03/Periodico_Salvador_Cumple.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.salvadorcumple.com/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2017/03/Periodico_Salvador_Cumple.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.salvadorcumple.com/#new_tab">Periódico Salvador Cumple</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2015/06/plan-quinquenal.jpg" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.presidencia.gob.sv/wp-content/uploads/2015/01/Plan-Quinquenal-de-Desarrollo.pdf#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2015/06/plan-quinquenal.jpg"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.presidencia.gob.sv/wp-content/uploads/2015/01/Plan-Quinquenal-de-Desarrollo.pdf#new_tab">Plan Quinquenal de Desarrollo 2014-2019</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2016/04/LOGO-PLAN-EL-SALVADOR-SEGURO.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://gobernabilidad.presidencia.gob.sv/plan-el-salvador-seguro/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2016/04/LOGO-PLAN-EL-SALVADOR-SEGURO.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://gobernabilidad.presidencia.gob.sv/plan-el-salvador-seguro/#new_tab">Plan El Salvador Seguro</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2014/12/Logo-GobSV.jpg" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://www.presidencia.gob.sv/directorio/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2014/12/Logo-GobSV.jpg"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://www.presidencia.gob.sv/directorio/#new_tab">Directorio Electrónico de Gobierno</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
									<li>
						<!-- THE MEDIA HOLDER PART -->
<div class="mediaholder">
	<div class="mediaholder_innerwrap">
		<img alt="image" src="http://www.salud.gob.sv/wp-content/uploads/2015/06/logo-canal-10-2016.png" style="height: auto;" width="290" height="155" >

		<!-- THE HOVER EFFECT (SPECIAL CLASS  - hovercover) -->
        <div class="hovercover">

			<!-- LINK TO THE POST -->
			<a href="http://tves.sv/#new_tab" target="_blank">
				<div class="linkicon notalone"><i class="sb-icon-link"></i></div>
			</a>
			<!-- LIGHTBOX LINK -->
			<a class="fancybox" rel="group" href="http://www.salud.gob.sv/wp-content/uploads/2015/06/logo-canal-10-2016.png"><div class="lupeicon notalone"><i class="sb-icon-search"></i></div></a>
		</div>	<!-- END OF THE HOVER EFFECT -->
      </div>
</div><!-- END OF MEDIA HOLDER PART -->

<!-- VISIBLE TEXTS ON THE TEASER - TITLE AND EXCERPT -->
<div class="detailholder">
	<div class="showbiz-title"><a href="http://tves.sv/#new_tab">Televisión de El Salvador</a></div>
	<div class="showbiz-description"></div>
</div>					</li>
					
				</ul>					
						<div class="sbclear"></div>
					</div> 
					<div class="sbclear"></div>
				</div>
				
									<!-- start navigation -->
					<div class="showbiz-navigation center">
	<a id="showbiz_left_1" class="sb-navigation-left"><i class="sb-icon-left-open"></i></a>
	<a id="showbiz_play_1" class="sb-navigation-play"><i class="sb-icon-play sb-playbutton"></i><i class="sb-icon-pause sb-pausebutton"></i></a>					
	<a id="showbiz_right_1" class="sb-navigation-right"><i class="sb-icon-right-open"></i></a>
	<div class="sbclear"></div>
</div>					<!--  end navigation -->
								
			</div>
			
						
						<script type="text/javascript">
			
							
				jQuery(document).ready(function() {
					
					if(jQuery('#showbiz_1_1').showbizpro == undefined)
						showbiz_showDoubleJqueryError('#showbiz_1_1');

					jQuery('#showbiz_1_1').showbizpro({
						dragAndScroll:"off",
						carousel:"on",
						allEntryAtOnce:"off",
						closeOtherOverlays:"off",
						entrySizeOffset:0,
						heightOffsetBottom:0,
						conteainerOffsetRight:0,
						forceFullWidth:false,
						visibleElementsArray:[4,3,2,1],
						rewindFromEnd:"off",
						autoPlay:"on",
						scrollOrientation:"left",						
						delay:"3000",
						speed:"300",
						easing:"Power1.easeOut"
					});
					
										
					jQuery(".fancybox").fancybox();
					
									});

			</script>
			
							
			<!-- END SHOWBIZ -->
			
			</div></div></div></div><div class="row vwpc-row"><div class="vwpc-section-custom_content"><div class="col-sm-12"><hr class="section-hr"><div class="pf-content"><div align="center">
<a href="https://www.facebook.com/ProgramaNacionaldeAlfabetizacionElSalvador/" target="_blank"><img src="/wp-content/uploads/2018/02/banner_ElSalvador-Alfabetizado.jpg" style="border: 1px solid #98181D; -webkit-border-radius: 10px; -moz-border-radius: 10px; border-radius: 10px; margin-bottom:10px;" title="El Salvador Alfabetizado | ¡es posible!"></a>
</div>
</div></div></div></div></div>

<hr>
<div class="col-sm-12" align="center">
<div align="center"><a href="http://www.isss.gob.sv/index.php?option=com_content&view=article&id=1608%25regimen-especial-para-salvadorenos-en-el-exterior&catid=103%25noticias-ciudadano&Itemid=77" target="_blank">
<img src="/wp-content/uploads/2017/12/Banner_ISSS_Regimen_Salud_503_1020x200.png" title="Régimen Salud 503 | Bienestar y tranquilidad para tu familia | Instituto Salvadoreño del Seguro Social ISSS"></a>
</div>
</div>
<hr>

<div class="col-sm-14" align="center">
<center>
<table border="0" cellspacing="0" cellpadding="0" width="100%" style="background-color:  #AEDEF1;">
  <tr>  
  <td align="center" valign="middle"><font color="#000000" face="Roboto" size="2">
   Contenido publicado bajo <a target=_new rel="license" href="http://creativecommons.org/licenses/by-sa/3.0/es/deed.es">licencia Creative Commons Atribución-CompartirIgual 3.0 Unported</a><br><img alt="Licencia Creative Commons" style="border-width:0" src="http://i.creativecommons.org/l/by-sa/3.0/80x15.png" /></a><br>(salvo donde específicamente se indiquen otros términos de licenciamiento)<br>
  Este sitio está totalmente basado en <a target=_new href="http://es.wikipedia.org/wiki/Software_libre"><b>Software Libre</b></a><br>[ <a target=_new href="http://www.debian.org">Debian GNU/Linux</a>, <a target=_new href="http://httpd.apache.org">Apache</a>, <a target=_new href="http://www.php.net">PHP</a>, <a target=_new href="http://www.mysql.com">MySQL</a> y <a target=_new href="https://es.wordpress.org/">Wordpress!</a> entre otros ]
</td>
</tr>
</table>
</center>
</div>				

<footer id="footer">
					<div class="footer-sidebar">
	<div class="container">
		<div class="row">
							<div class="footer-sidebar-1 widget-area col-sm-4" role="complementary">
				<div id="custom_html-6" class="widget_text widget vw-sidebar-footer-1 widget_custom_html"><div class="textwidget custom-html-widget"><div align="center">
<a href="http://www.presidencia.gob.sv" target="_blank"><img src="/images/escudo-el-salvador-oficial-peque.png" alt="Presidencia de la República" title="Presidencia de la República de El Salvador"></a></div></div></div>				</div>
			
							<div class="footer-sidebar-2 widget-area col-sm-4" role="complementary">
				<div id="custom_html-7" class="widget_text widget vw-sidebar-footer-2 widget_custom_html"><div class="textwidget custom-html-widget"><div align="center">
<b>Ministerio de Salud<br>
REPÚBLICA DE EL SALVADOR, C.A.<br>
Calle Arce No.827, San Salvador, El Salvador, C.A.<br>
Conmutador: (503) 2591-7000 • Fax: (503) 2221-0991.</b>
</div>

<div align="center"><font face="Verdana" size="1">
<img src="/images/email_white.png" title="Contáctenos">&nbsp;<a href="/contactenos-unidad-por-el-derecho-a-la-salud/" title="Contáctenos">Contáctenos</a> | <img src="/images/email_white.png" title="Webmaster">&nbsp;<a href="/webmaster/" title="Webmaster">Webmaster</a><br><a href="/politica-web/" title="Política de Seguridad y Privacidad del MINSAL - El Salvador">Política de Seguridad y Privacidad</a></font>
</div></div></div>				</div>
			
							<div class="footer-sidebar-3 widget-area col-sm-4" role="complementary">
				<div id="custom_html-8" class="widget_text widget vw-sidebar-footer-3 widget_custom_html"><div class="textwidget custom-html-widget"><div align="center"><a rel="nofollow" title="Estandarización de Sitios Web" href="http://estandarizacion.itiges.sv/?p=332" target="_blank"><img alt="Estandarización de Sitios Web" src="/images/boton_estandarizado2.0_minsal.png" ></a>
</div></div></div>				</div>
					</div>
	</div>
</div>

					<div class="copyright">
						<div class="container">
							<div class="row">
								<div class="col-sm-6 copyright-left"><a href="/derechos-de-informacion/">Derechos de Información 2017.</a> Ministerio de Salud de El Salvador.</div>
								<div class="col-sm-6 copyright-right">
									<a class="back-to-top" href="#top">&uarr;	Subir</a>
								</div>
							</div>
						</div>
					</div>
				</footer>
			
			</div> <!-- Off canvas body inner -->
		<script type="text/html" id="tmpl-wp-playlist-current-item">
	<# if ( data.image ) { #>
	<img src="{{ data.thumb.src }}" alt="" />
	<# } #>
	<div class="wp-playlist-caption">
		<span class="wp-playlist-item-meta wp-playlist-item-title">&#8220;{{ data.title }}&#8221;</span>
		<# if ( data.meta.album ) { #><span class="wp-playlist-item-meta wp-playlist-item-album">{{ data.meta.album }}</span><# } #>
		<# if ( data.meta.artist ) { #><span class="wp-playlist-item-meta wp-playlist-item-artist">{{ data.meta.artist }}</span><# } #>
	</div>
</script>
<script type="text/html" id="tmpl-wp-playlist-item">
	<div class="wp-playlist-item">
		<a class="wp-playlist-caption" href="{{ data.src }}">
			{{ data.index ? ( data.index + '. ' ) : '' }}
			<# if ( data.caption ) { #>
				{{ data.caption }}
			<# } else { #>
				<span class="wp-playlist-item-title">&#8220;{{{ data.title }}}&#8221;</span>
				<# if ( data.artists && data.meta.artist ) { #>
				<span class="wp-playlist-item-artist"> &mdash; {{ data.meta.artist }}</span>
				<# } #>
			<# } #>
		</a>
		<# if ( data.meta.length_formatted ) { #>
		<div class="wp-playlist-item-length">{{ data.meta.length_formatted }}</div>
		<# } #>
	</div>
</script>
<script type="text/javascript">

  var _gaq = _gaq || [];
  _gaq.push(['_setAccount', 'UA-20729832-1']);
  _gaq.push(['_trackPageview']);

  (function() {
    var ga = document.createElement('script'); ga.type = 'text/javascript'; ga.async = true;
    ga.src = ('https:' == document.location.protocol ? 'https://ssl' : 'http://www') + '.google-analytics.com/ga.js';
    var s = document.getElementsByTagName('script')[0]; s.parentNode.insertBefore(ga, s);
  })();

</script>		<script type='text/javascript'>
			;(function( $, window, document, undefined ){
				"use strict";

				$( document ).ready( function ($) {
							$( '.flexslider' ).flexslider({
			animation: "fade",
			easing: "easeInCirc",
			slideshow: true,
			slideshowSpeed: 4000,
			animationSpeed: 600,
			randomize: false,
			pauseOnHover: true,
			prevText: '',
			nextText: '',
			start: function( slider ) {
				slider.css( 'opacity', '1' );
				slider.find( '.post-thumbnail-wrapper' ).css( 'height', '500px' ).imgLiquid().fadeIn(250);
			},
		});
					} );
				
			})( jQuery, window , document );

					</script>
		    <script>jQuery(document).ready(function($) { $('#flags a, a.single-language, .tool-items a').each(function() { $(this).attr('data-lang', $(this).attr('title')); }); $(document.body).on("click","a.flag", function(){function l(){doGoogleLanguageTranslator(default_lang+"|"+default_lang); }function n(){doGoogleLanguageTranslator(default_lang+"|"+lang_prefix); } lang_text=$(this).attr('data-lang'),default_lang="es",lang_prefix=$(this).attr("class").split(" ")[2],$(".tool-container").hide(),lang_prefix==default_lang?l():n()}),0==$("body > #google_language_translator").length&&$("#glt-footer").html("<div id='google_language_translator'></div>"); });</script><script type='text/javascript' src='//translate.google.com/translate_a/element.js?cb=GoogleLanguageTranslatorInit'></script>

    <div id="flags" style="display:none" class="size18"><ul id="sortable" class="ui-sortable"></ul></div><div id='glt-footer'></div><script type='text/javascript'>function GoogleLanguageTranslatorInit() { new google.translate.TranslateElement({pageLanguage: 'es', includedLanguages:'af,sq,am,ar,hy,az,eu,be,bn,bs,bg,ca,ceb,ny,zh-CN,zh-TW,co,hr,cs,da,nl,en,eo,et,tl,fi,fr,fy,gl,ka,de,el,gu,ht,ha,haw,iw,hi,hmn,hu,is,ig,id,ga,it,ja,jw,kn,kk,km,ko,ku,ky,lo,la,lv,lt,lb,mk,mg,ml,ms,mt,mi,mr,mn,my,ne,no,ps,fa,pl,pt,pa,ro,ru,sr,sn,st,sd,si,sk,sl,sm,gd,so,es,su,sw,sv,tg,ta,te,th,tr,uk,ur,uz,vi,cy,xh,yi,yo,zu', autoDisplay: false, multilanguagePage:true}, 'google_language_translator');}</script><div class="scroll-back-to-top-wrapper">
	<span class="scroll-back-to-top-inner">
					<i class="fa fa-2x fa-arrow-circle-up"></i>
			</span>
</div>        <div class="w3eden">
            <div id="wpdm-popup-link" class="modal fade">
                <div class="modal-dialog" style="width: 750px">
                    <div class="modal-content">
                        <div class="modal-header">
                              <h4 class="modal-title"></h4>
                        </div>
                        <div class="modal-body" id='wpdm-modal-body'>
                            <p class="placeholder">
                                [ Placeholder content for popup link ]
                                <a href="https://www.wpdownloadmanager.com/">WordPress Download Manager - Best Download Management Plugin</a>
                            </p>
                        </div>
                        <div class="modal-footer">
                            <button type="button" class="btn btn-danger" data-dismiss="modal">Close</button>
                        </div>
                    </div><!-- /.modal-content -->
                </div><!-- /.modal-dialog -->
            </div><!-- /.modal -->


        </div>
        <script language="JavaScript">
            <!--
            jQuery(function () {
                jQuery('.wpdm-popup-link').click(function (e) {
                    e.preventDefault();
                    jQuery('#wpdm-popup-link .modal-title').html(jQuery(this).data('title'));
                    jQuery('#wpdm-modal-body').html('<i class="icon"><img align="left" style="margin-top: -1px" src="http://www.salud.gob.sv/wp-content/plugins/download-manager/assets/images/loading-new.gif" /></i>&nbsp;Please Wait...');
                    jQuery('#wpdm-popup-link').modal('show');
                    jQuery.post(this.href,{mode:'popup'}, function (res) {
                        jQuery('#wpdm-modal-body').html(res);
                    });
                    return false;
                });
            });
            //-->
        </script>
        <style type="text/css">
            #wpdm-modal-body img {
                max-width: 100% !important;
            }
            .placeholder{
                display: none;
            }
        </style>
    		<script>
		( function ( body ) {
			'use strict';
			body.className = body.className.replace( /\btribe-no-js\b/, 'tribe-js' );
		} )( document.body );
		</script>
		<script type='text/javascript'> /* <![CDATA[ */var tribe_l10n_datatables = {"aria":{"sort_ascending":": activate to sort column ascending","sort_descending":": activate to sort column descending"},"length_menu":"Show _MENU_ entries","empty_table":"No data available in table","info":"Showing _START_ to _END_ of _TOTAL_ entries","info_empty":"Showing 0 to 0 of 0 entries","info_filtered":"(filtered from _MAX_ total entries)","zero_records":"No matching records found","search":"Search:","all_selected_text":"All items on this page were selected. ","select_all_link":"Select all pages","clear_selection":"Clear Selection.","pagination":{"all":"All","next":"Next","previous":"Previous"},"select":{"rows":{"0":"","_":": Selected %d rows","1":": Selected 1 row"}},"datepicker":{"dayNames":["domingo","lunes","martes","mi\u00e9rcoles","jueves","viernes","s\u00e1bado"],"dayNamesShort":["Dom","Lun","Mar","Mie","Jue","Vie","Sab"],"dayNamesMin":["D","L","M","X","J","V","S"],"monthNames":["enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre"],"monthNamesShort":["enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre"],"nextText":"Siguiente","prevText":"Anterior","currentText":"Hoy","closeText":"Hecho"}};/* ]]> */ </script>      <script type="text/javascript">

          var pfHeaderImgUrl = '';
          var pfHeaderTagline = '';
          var pfdisableClickToDel = '1';
          var pfImagesSize = 'full-size';
          var pfImageDisplayStyle = 'block';
          var pfDisableEmail = '0';
          var pfDisablePDF = '0';
          var pfDisablePrint = '0';
          var pfCustomCSS = '';
          var pfPlatform = 'Wordpress';
      (function() {
            var e = document.createElement('script'); e.type="text/javascript";
            e.src = 'https://cdn.printfriendly.com/printfriendly.js';
            document.getElementsByTagName('head')[0].appendChild(e);
        })();
      </script>
<link rel='stylesheet' id='mediaelement-css'  href='http://www.salud.gob.sv/wp-includes/js/mediaelement/mediaelementplayer-legacy.min.css?ver=4.2.6-78496d1' type='text/css' media='all' />
<link rel='stylesheet' id='wp-mediaelement-css'  href='http://www.salud.gob.sv/wp-includes/js/mediaelement/wp-mediaelement.min.css?ver=4.9.4' type='text/css' media='all' />
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/comment-reply.min.js?ver=4.9.4'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var wpcf7 = {"apiSettings":{"root":"http:\/\/www.salud.gob.sv\/wp-json\/contact-form-7\/v1","namespace":"contact-form-7\/v1"},"recaptcha":{"messages":{"empty":"Por favor, prueba que no eres un robot."}},"cached":"1"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/contact-form-7/includes/js/scripts.js?ver=5.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/core.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/datepicker.min.js?ver=1.11.4'></script>
<script type='text/javascript'>
jQuery(document).ready(function(jQuery){jQuery.datepicker.setDefaults({"closeText":"Cerrar","currentText":"Hoy","monthNames":["enero","febrero","marzo","abril","mayo","junio","julio","agosto","septiembre","octubre","noviembre","diciembre"],"monthNamesShort":["Ene","Feb","Mar","Abr","May","Jun","Jul","Ago","Sep","Oct","Nov","Dic"],"nextText":"Siguiente","prevText":"Previo","dayNames":["domingo","lunes","martes","mi\u00e9rcoles","jueves","viernes","s\u00e1bado"],"dayNamesShort":["Dom","Lun","Mar","Mie","Jue","Vie","Sab"],"dayNamesMin":["D","L","M","X","J","V","S"],"dateFormat":"d MM, yy","firstDay":1,"isRTL":false});});
</script>
<script type='text/javascript' src='http://ajax.googleapis.com/ajax/libs/jqueryui/1.11.4/i18n/datepicker-es.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/contact-form-7-datepicker/js/jquery-ui-timepicker/jquery-ui-timepicker-addon.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/contact-form-7-datepicker/js/jquery-ui-timepicker/i18n/jquery-ui-timepicker-es.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/widget.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/mouse.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/slider.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/button.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/contact-form-7-datepicker/js/jquery-ui-sliderAccess.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/jquery.form.min.js?ver=4.2.1'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var scrollBackToTop = {"scrollDuration":"500","fadeDuration":"0.5"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/scroll-back-to-top/assets/js/scroll-back-to-top.js'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/zeno-font-resizer/js/js.cookie.js?ver=1.7.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/zeno-font-resizer/js/jquery.fontsize.js?ver=1.7.1'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var spuvar = {"is_admin":"","disable_style":"","safe_mode":"","ajax_mode":"","ajax_url":"http:\/\/www.salud.gob.sv\/wp-admin\/admin-ajax.php","ajax_mode_url":"http:\/\/www.salud.gob.sv\/?spu_action=spu_load&lang=","pid":"15","is_front_page":"1","is_category":"","site_url":"http:\/\/www.salud.gob.sv","is_archive":"","is_search":"","is_preview":"","seconds_confirmation_close":"5"};
var spuvar_social = [];
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/popups/public/assets/js/min/public-min.js?ver=1.9.1.1'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var pplb_ajax = {"ajaxurl":"http:\/\/www.salud.gob.sv\/wp-admin\/admin-ajax.php"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/protected-posts-logout-button/logout.js'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/page-links-to/js/new-tab.min.js?ver=2.9.8'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/effect.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/jquery/ui/effect-fade.min.js?ver=1.11.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/js/jquery.fitvids.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/js/jquery.isotope.min.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/flexslider/jquery.flexslider.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/framework/swipebox/jquery.swipebox.min.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/js/asset.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/themes/RedSV/js/main.js?ver=1.9.0'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/js/bootstrap-dropdown.js?ver=3.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/js/bootstrap-tab.js?ver=3.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/js/bootstrap-tabdrop.js?ver=3.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/easy-responsive-tabs/assets/js/ert_js.php?ver=3.1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/hoverIntent.min.js?ver=1.8.1'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var megamenu = {"timeout":"300","interval":"100"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/megamenu/js/maxmegamenu.js?ver=2.4.1.2'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/wp-embed.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-content/plugins/the-events-calendar/common/src/resources/js/underscore-before.js'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/underscore.min.js?ver=1.8.3'></script>
<script type='text/Javascript' src='http://www.salud.gob.sv/wp-content/plugins/the-events-calendar/common/src/resources/js/underscore-after.js'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var _wpUtilSettings = {"ajax":{"url":"\/wp-admin\/admin-ajax.php"}};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/wp-util.min.js?ver=4.9.4'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/backbone.min.js?ver=1.2.3'></script>
<script type='text/javascript'>
var mejsL10n = {"language":"es","strings":{"mejs.install-flash":"Est\u00e1s usando un navegador que no tiene Flash activo o instalado. Por favor, activa el componente del reproductor Flash o descarga la \u00faltima versi\u00f3n desde https:\/\/get.adobe.com\/flashplayer\/","mejs.fullscreen-off":"Salir de pantalla completa","mejs.fullscreen-on":"Ver en pantalla completa","mejs.download-video":"Descargar v\u00eddeo","mejs.fullscreen":"Pantalla completa","mejs.time-jump-forward":["Saltar %1 segundo hacia adelante","Salta hacia adelante %1 segundos"],"mejs.loop":"Alternar bucle","mejs.play":"Reproducir","mejs.pause":"Pausa","mejs.close":"Cerrar","mejs.time-slider":"Control de tiempo","mejs.time-help-text":"Usa las teclas de direcci\u00f3n izquierda\/derecha para avanzar un segundo, y las flechas arriba\/abajo para avanzar diez segundos.","mejs.time-skip-back":["Saltar atr\u00e1s 1 segundo","Retroceder %1 segundos"],"mejs.captions-subtitles":"Pies de foto \/ Subt\u00edtulos","mejs.captions-chapters":"Cap\u00edtulos","mejs.none":"Ninguna","mejs.mute-toggle":"Desactivar sonido","mejs.volume-help-text":"Utiliza las teclas de flecha arriba\/abajo para aumentar o disminuir el volumen.","mejs.unmute":"Activar sonido","mejs.mute":"Silenciar","mejs.volume-slider":"Control de volumen","mejs.video-player":"Reproductor de v\u00eddeo","mejs.audio-player":"Reproductor de audio","mejs.ad-skip":"Saltar anuncio","mejs.ad-skip-info":["Saltar en 1 segundo","Saltar en %1 segundos"],"mejs.source-chooser":"Selector de origen","mejs.stop":"Parar","mejs.speed-rate":"Tasa de velocidad","mejs.live-broadcast":"Transmisi\u00f3n en vivo","mejs.afrikaans":"Africano","mejs.albanian":"Albano","mejs.arabic":"\u00c1rabe","mejs.belarusian":"Bielorruso","mejs.bulgarian":"B\u00falgaro","mejs.catalan":"Catal\u00e1n","mejs.chinese":"Chino","mejs.chinese-simplified":"Chino (Simplificado)","mejs.chinese-traditional":"Chino (Tradicional)","mejs.croatian":"Croata","mejs.czech":"Checo","mejs.danish":"Dan\u00e9s","mejs.dutch":"Holand\u00e9s","mejs.english":"Ingl\u00e9s","mejs.estonian":"Estonio","mejs.filipino":"Filipino","mejs.finnish":"Fin\u00e9s","mejs.french":"Franc\u00e9s","mejs.galician":"Gallego","mejs.german":"Alem\u00e1n","mejs.greek":"Griego","mejs.haitian-creole":"Creole haitiano","mejs.hebrew":"Hebreo","mejs.hindi":"Indio","mejs.hungarian":"H\u00fangaro","mejs.icelandic":"Island\u00e9s","mejs.indonesian":"Indonesio","mejs.irish":"Irland\u00e9s","mejs.italian":"Italiano","mejs.japanese":"Japon\u00e9s","mejs.korean":"Coreano","mejs.latvian":"Let\u00f3n","mejs.lithuanian":"Lituano","mejs.macedonian":"Macedonio","mejs.malay":"Malayo","mejs.maltese":"Malt\u00e9s","mejs.norwegian":"Noruego","mejs.persian":"Persa","mejs.polish":"Polaco","mejs.portuguese":"Portugu\u00e9s","mejs.romanian":"Rumano","mejs.russian":"Ruso","mejs.serbian":"Serbio","mejs.slovak":"Eslovaco","mejs.slovenian":"Esloveno","mejs.spanish":"Espa\u00f1ol","mejs.swahili":"Swahili","mejs.swedish":"Sueco","mejs.tagalog":"Tagalo","mejs.thai":"Thai","mejs.turkish":"Turco","mejs.ukrainian":"Ukraniano","mejs.vietnamese":"Vietnamita","mejs.welsh":"Gal\u00e9s","mejs.yiddish":"Yiddish"}};
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/mediaelement/mediaelement-and-player.min.js?ver=4.2.6-78496d1'></script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/mediaelement/mediaelement-migrate.min.js?ver=4.9.4'></script>
<script type='text/javascript'>
/* <![CDATA[ */
var _wpmejsSettings = {"pluginPath":"\/wp-includes\/js\/mediaelement\/","classPrefix":"mejs-","stretching":"responsive"};
/* ]]> */
</script>
<script type='text/javascript' src='http://www.salud.gob.sv/wp-includes/js/mediaelement/wp-playlist.min.js?ver=4.9.4'></script>
	</body>
</html>